/*
    Shama v1.0.0, for tinytapeout3.
    Copyright (C) 2023 Pat Deegan, https://psychogenic.com
    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.
    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.
    You should have received a copy of the GNU General Public License
    along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/

`default_nettype none
`timescale 1ns/1ps
/* Generated by Amaranth Yosys 0.25 (PyPI ver 0.25.0.0.post69, git sha1 e02b7f64b) */

module \buf ();
  wire \$empty_module_filler ;
endmodule

module ch(ch_y, ch_z, ch_out, ch_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  wire [31:0] \$7 ;
  output [31:0] ch_out;
  wire [31:0] ch_out;
  input [31:0] ch_x;
  wire [31:0] ch_x;
  input [31:0] ch_y;
  wire [31:0] ch_y;
  input [31:0] ch_z;
  wire [31:0] ch_z;
  assign \$1  = ch_x & ch_y;
  assign \$3  = ~ ch_x;
  assign \$5  = \$3  & ch_z;
  assign \$7  = \$1  ^ \$5 ;
  assign ch_out = \$7 ;
endmodule

module maj(maj_y, maj_z, maj_out, maj_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  wire [31:0] \$7 ;
  wire [31:0] \$9 ;
  output [31:0] maj_out;
  wire [31:0] maj_out;
  input [31:0] maj_x;
  wire [31:0] maj_x;
  input [31:0] maj_y;
  wire [31:0] maj_y;
  input [31:0] maj_z;
  wire [31:0] maj_z;
  assign \$9  = \$5  ^ \$7 ;
  assign \$1  = maj_x & maj_y;
  assign \$3  = maj_x & maj_z;
  assign \$5  = \$1  ^ \$3 ;
  assign \$7  = maj_y & maj_z;
  assign maj_out = \$9 ;
endmodule

module nibbler(rst, inNibble, inputReady, busy, nres_out, clk);
  reg \$auto$verilog_backend.cc:2083:dump_module$1  = 0;
  wire [34:0] \$1 ;
  wire [34:0] \$10 ;
  wire \$1000 ;
  wire \$1002 ;
  wire \$1004 ;
  wire \$1006 ;
  wire [9:0] \$1008 ;
  wire [9:0] \$1009 ;
  wire \$101 ;
  wire \$1011 ;
  wire \$1013 ;
  wire \$1015 ;
  wire \$1017 ;
  wire \$1019 ;
  wire \$1021 ;
  wire \$1023 ;
  wire \$1025 ;
  wire \$1027 ;
  wire \$1029 ;
  wire \$103 ;
  wire \$1031 ;
  wire \$1033 ;
  wire \$1035 ;
  wire \$1037 ;
  wire \$1039 ;
  wire \$1041 ;
  wire \$1043 ;
  wire \$1045 ;
  wire \$1047 ;
  wire \$1049 ;
  wire \$105 ;
  wire \$1051 ;
  wire \$1053 ;
  wire \$1055 ;
  wire \$1057 ;
  wire \$1059 ;
  wire \$1061 ;
  wire \$1063 ;
  wire \$1065 ;
  wire \$1067 ;
  wire \$1069 ;
  wire \$107 ;
  wire \$1071 ;
  wire \$1073 ;
  wire \$1075 ;
  wire \$1077 ;
  wire \$1079 ;
  wire \$1081 ;
  wire \$1083 ;
  wire \$1085 ;
  wire \$1087 ;
  wire \$1089 ;
  wire \$109 ;
  wire \$1091 ;
  wire \$1093 ;
  wire \$1095 ;
  wire \$1097 ;
  wire \$1099 ;
  wire \$1101 ;
  wire \$1103 ;
  wire \$1105 ;
  wire \$1107 ;
  wire \$1109 ;
  wire \$111 ;
  wire \$1111 ;
  wire \$1113 ;
  wire \$1115 ;
  wire \$1117 ;
  wire \$1119 ;
  wire \$1121 ;
  wire \$1123 ;
  wire \$1125 ;
  wire \$1127 ;
  wire \$1129 ;
  wire \$113 ;
  wire \$1131 ;
  wire \$1133 ;
  wire \$1135 ;
  wire \$1137 ;
  wire [32:0] \$1139 ;
  wire [32:0] \$1140 ;
  wire \$1142 ;
  wire \$1144 ;
  wire \$1146 ;
  wire \$1148 ;
  wire \$115 ;
  wire \$1150 ;
  wire \$1152 ;
  wire \$117 ;
  wire \$119 ;
  wire [34:0] \$12 ;
  wire \$121 ;
  wire \$123 ;
  wire \$125 ;
  wire \$127 ;
  wire \$129 ;
  wire \$131 ;
  wire \$133 ;
  wire \$135 ;
  wire \$137 ;
  wire \$139 ;
  wire [34:0] \$14 ;
  wire \$141 ;
  wire \$143 ;
  wire \$145 ;
  wire \$147 ;
  wire \$149 ;
  wire \$151 ;
  wire \$153 ;
  wire \$155 ;
  wire \$157 ;
  wire \$159 ;
  wire [18:0] \$16 ;
  wire \$161 ;
  wire \$163 ;
  wire \$165 ;
  wire [31:0] \$167 ;
  wire [31:0] \$168 ;
  wire [31:0] \$170 ;
  wire \$172 ;
  wire [31:0] \$174 ;
  wire [31:0] \$175 ;
  wire [31:0] \$177 ;
  wire \$179 ;
  wire [34:0] \$18 ;
  wire [31:0] \$181 ;
  wire [31:0] \$182 ;
  wire [31:0] \$184 ;
  wire \$186 ;
  wire [31:0] \$188 ;
  wire [31:0] \$189 ;
  wire [31:0] \$191 ;
  wire \$193 ;
  wire [31:0] \$195 ;
  wire [31:0] \$196 ;
  wire [31:0] \$198 ;
  wire [34:0] \$2 ;
  wire [18:0] \$20 ;
  wire \$200 ;
  wire [31:0] \$202 ;
  wire [31:0] \$203 ;
  wire [31:0] \$205 ;
  wire \$207 ;
  wire [31:0] \$209 ;
  wire [31:0] \$210 ;
  wire [31:0] \$212 ;
  wire \$214 ;
  wire [31:0] \$216 ;
  wire [31:0] \$217 ;
  wire [31:0] \$219 ;
  wire [34:0] \$22 ;
  wire \$221 ;
  wire [31:0] \$223 ;
  wire [31:0] \$224 ;
  wire [31:0] \$226 ;
  wire \$228 ;
  wire [31:0] \$230 ;
  wire [31:0] \$231 ;
  wire [31:0] \$233 ;
  wire \$235 ;
  wire [31:0] \$237 ;
  wire [31:0] \$238 ;
  wire [10:0] \$24 ;
  wire [31:0] \$240 ;
  wire \$242 ;
  wire [31:0] \$244 ;
  wire [31:0] \$245 ;
  wire [31:0] \$247 ;
  wire \$249 ;
  wire [31:0] \$251 ;
  wire [31:0] \$252 ;
  wire [31:0] \$254 ;
  wire \$256 ;
  wire [31:0] \$258 ;
  wire [31:0] \$259 ;
  wire [34:0] \$26 ;
  wire [31:0] \$261 ;
  wire \$263 ;
  wire [31:0] \$265 ;
  wire [31:0] \$266 ;
  wire [31:0] \$268 ;
  wire \$270 ;
  wire [31:0] \$272 ;
  wire [31:0] \$273 ;
  wire [31:0] \$275 ;
  wire \$277 ;
  wire [31:0] \$279 ;
  wire [34:0] \$28 ;
  wire [31:0] \$280 ;
  wire [31:0] \$282 ;
  wire \$284 ;
  wire [31:0] \$286 ;
  wire [31:0] \$287 ;
  wire [31:0] \$289 ;
  wire \$291 ;
  wire [31:0] \$293 ;
  wire [31:0] \$294 ;
  wire [31:0] \$296 ;
  wire \$298 ;
  wire [6:0] \$30 ;
  wire [31:0] \$300 ;
  wire [31:0] \$301 ;
  wire [31:0] \$303 ;
  wire \$305 ;
  wire [31:0] \$307 ;
  wire [31:0] \$308 ;
  wire [6:0] \$31 ;
  wire [31:0] \$310 ;
  wire \$312 ;
  wire [31:0] \$314 ;
  wire [31:0] \$315 ;
  wire [31:0] \$317 ;
  wire \$319 ;
  wire [31:0] \$321 ;
  wire [31:0] \$322 ;
  wire [31:0] \$324 ;
  wire \$326 ;
  wire [31:0] \$328 ;
  wire [31:0] \$329 ;
  wire \$33 ;
  wire [31:0] \$331 ;
  wire \$333 ;
  wire [31:0] \$335 ;
  wire [31:0] \$336 ;
  wire [31:0] \$338 ;
  wire \$340 ;
  wire [31:0] \$342 ;
  wire [31:0] \$343 ;
  wire [31:0] \$345 ;
  wire \$347 ;
  wire [31:0] \$349 ;
  wire \$35 ;
  wire [31:0] \$350 ;
  wire [31:0] \$352 ;
  wire \$354 ;
  wire [31:0] \$356 ;
  wire [31:0] \$357 ;
  wire [31:0] \$359 ;
  wire \$361 ;
  wire [31:0] \$363 ;
  wire [31:0] \$364 ;
  wire [31:0] \$366 ;
  wire \$368 ;
  wire \$37 ;
  wire [31:0] \$370 ;
  wire [31:0] \$371 ;
  wire [31:0] \$373 ;
  wire \$375 ;
  wire [31:0] \$377 ;
  wire [31:0] \$378 ;
  wire [31:0] \$380 ;
  wire \$382 ;
  wire [31:0] \$384 ;
  wire [31:0] \$385 ;
  wire [31:0] \$387 ;
  wire \$389 ;
  wire \$39 ;
  wire [31:0] \$391 ;
  wire [31:0] \$392 ;
  wire [31:0] \$394 ;
  wire \$396 ;
  wire [31:0] \$398 ;
  wire [31:0] \$399 ;
  wire [34:0] \$4 ;
  wire [31:0] \$401 ;
  wire \$403 ;
  wire [31:0] \$405 ;
  wire [31:0] \$406 ;
  wire [31:0] \$408 ;
  wire \$41 ;
  wire \$410 ;
  wire [31:0] \$412 ;
  wire [31:0] \$413 ;
  wire [31:0] \$415 ;
  wire \$417 ;
  wire [31:0] \$419 ;
  wire [31:0] \$420 ;
  wire [31:0] \$422 ;
  wire \$424 ;
  wire [31:0] \$426 ;
  wire [31:0] \$427 ;
  wire [31:0] \$429 ;
  wire \$43 ;
  wire \$431 ;
  wire [31:0] \$433 ;
  wire [31:0] \$434 ;
  wire [31:0] \$436 ;
  wire \$438 ;
  wire [31:0] \$440 ;
  wire [31:0] \$441 ;
  wire [31:0] \$443 ;
  wire \$445 ;
  wire [31:0] \$447 ;
  wire [31:0] \$448 ;
  wire \$45 ;
  wire [31:0] \$450 ;
  wire \$452 ;
  wire [31:0] \$454 ;
  wire [31:0] \$455 ;
  wire [31:0] \$457 ;
  wire \$459 ;
  wire [31:0] \$461 ;
  wire [31:0] \$462 ;
  wire [31:0] \$464 ;
  wire \$466 ;
  wire [31:0] \$468 ;
  wire [31:0] \$469 ;
  wire \$47 ;
  wire [31:0] \$471 ;
  wire \$473 ;
  wire [31:0] \$475 ;
  wire [31:0] \$476 ;
  wire [31:0] \$478 ;
  wire \$480 ;
  wire [31:0] \$482 ;
  wire [31:0] \$483 ;
  wire [31:0] \$485 ;
  wire \$487 ;
  wire [31:0] \$489 ;
  wire \$49 ;
  wire [31:0] \$490 ;
  wire [31:0] \$492 ;
  wire \$494 ;
  wire [31:0] \$496 ;
  wire [31:0] \$497 ;
  wire [31:0] \$499 ;
  wire \$501 ;
  wire [31:0] \$503 ;
  wire [31:0] \$504 ;
  wire [31:0] \$506 ;
  wire \$508 ;
  wire \$51 ;
  wire [31:0] \$510 ;
  wire [31:0] \$511 ;
  wire [31:0] \$513 ;
  wire \$515 ;
  wire [31:0] \$517 ;
  wire [31:0] \$518 ;
  wire [31:0] \$520 ;
  wire \$522 ;
  wire [31:0] \$524 ;
  wire [31:0] \$525 ;
  wire [31:0] \$527 ;
  wire \$529 ;
  wire \$53 ;
  wire [31:0] \$531 ;
  wire [31:0] \$532 ;
  wire [31:0] \$534 ;
  wire \$536 ;
  wire [31:0] \$538 ;
  wire [31:0] \$539 ;
  wire [31:0] \$541 ;
  wire \$543 ;
  wire [31:0] \$545 ;
  wire [31:0] \$546 ;
  wire [31:0] \$548 ;
  wire \$55 ;
  wire \$550 ;
  wire [31:0] \$552 ;
  wire [31:0] \$553 ;
  wire [31:0] \$555 ;
  wire \$557 ;
  wire [31:0] \$559 ;
  wire [31:0] \$560 ;
  wire [31:0] \$562 ;
  wire \$564 ;
  wire [31:0] \$566 ;
  wire [31:0] \$567 ;
  wire [31:0] \$569 ;
  wire \$57 ;
  wire \$571 ;
  wire [31:0] \$573 ;
  wire [31:0] \$574 ;
  wire [31:0] \$576 ;
  wire \$578 ;
  wire [31:0] \$580 ;
  wire [31:0] \$581 ;
  wire [31:0] \$583 ;
  wire \$585 ;
  wire [31:0] \$587 ;
  wire [31:0] \$588 ;
  wire \$59 ;
  wire [31:0] \$590 ;
  wire \$592 ;
  wire [31:0] \$594 ;
  wire [31:0] \$595 ;
  wire [31:0] \$597 ;
  wire \$599 ;
  wire [34:0] \$6 ;
  wire [31:0] \$601 ;
  wire [31:0] \$602 ;
  wire [31:0] \$604 ;
  wire \$606 ;
  wire [31:0] \$608 ;
  wire [31:0] \$609 ;
  wire \$61 ;
  wire [31:0] \$611 ;
  wire \$613 ;
  wire \$615 ;
  wire \$617 ;
  wire \$619 ;
  wire \$621 ;
  wire \$623 ;
  wire \$625 ;
  wire \$627 ;
  wire \$629 ;
  wire \$63 ;
  wire \$631 ;
  wire \$633 ;
  wire \$635 ;
  wire \$637 ;
  wire \$639 ;
  wire \$641 ;
  wire \$643 ;
  wire \$645 ;
  wire \$647 ;
  wire \$649 ;
  wire \$65 ;
  wire \$651 ;
  wire \$653 ;
  wire \$655 ;
  wire \$657 ;
  wire \$659 ;
  wire \$661 ;
  wire \$663 ;
  wire \$665 ;
  wire \$667 ;
  wire [4:0] \$669 ;
  wire \$67 ;
  wire [4:0] \$670 ;
  wire \$672 ;
  wire \$674 ;
  wire \$676 ;
  wire [8:0] \$678 ;
  wire [8:0] \$679 ;
  wire \$681 ;
  wire \$683 ;
  wire \$685 ;
  wire \$687 ;
  wire \$689 ;
  wire \$69 ;
  wire \$691 ;
  wire \$693 ;
  wire \$695 ;
  wire \$697 ;
  wire \$699 ;
  wire \$701 ;
  wire \$703 ;
  wire \$705 ;
  wire \$707 ;
  wire \$709 ;
  wire \$71 ;
  wire \$711 ;
  wire \$713 ;
  wire \$715 ;
  wire \$717 ;
  wire \$719 ;
  wire \$721 ;
  wire \$723 ;
  wire [574:0] \$725 ;
  wire [574:0] \$726 ;
  wire [574:0] \$728 ;
  wire \$73 ;
  wire \$730 ;
  wire \$732 ;
  wire [5:0] \$734 ;
  wire [5:0] \$735 ;
  wire \$737 ;
  wire [7:0] \$739 ;
  wire [7:0] \$740 ;
  wire [32:0] \$742 ;
  wire [32:0] \$743 ;
  wire [32:0] \$745 ;
  wire [32:0] \$746 ;
  wire [32:0] \$748 ;
  wire [32:0] \$749 ;
  wire \$75 ;
  wire [32:0] \$751 ;
  wire [32:0] \$752 ;
  wire [32:0] \$754 ;
  wire [32:0] \$755 ;
  wire [32:0] \$757 ;
  wire [32:0] \$758 ;
  wire [32:0] \$760 ;
  wire [32:0] \$761 ;
  wire [32:0] \$763 ;
  wire [32:0] \$764 ;
  wire \$766 ;
  wire \$768 ;
  wire \$77 ;
  wire [32:0] \$770 ;
  wire [32:0] \$771 ;
  wire [32:0] \$773 ;
  wire [32:0] \$774 ;
  wire \$776 ;
  wire \$778 ;
  wire [4:0] \$780 ;
  wire [4:0] \$781 ;
  wire \$783 ;
  wire \$785 ;
  wire [35:0] \$787 ;
  wire [32:0] \$788 ;
  wire \$79 ;
  wire [33:0] \$790 ;
  wire [34:0] \$792 ;
  wire [35:0] \$794 ;
  wire \$796 ;
  wire \$798 ;
  wire [34:0] \$8 ;
  wire \$800 ;
  wire \$802 ;
  wire \$804 ;
  wire \$806 ;
  wire \$808 ;
  wire \$81 ;
  wire \$810 ;
  wire \$812 ;
  wire \$814 ;
  wire \$816 ;
  wire \$818 ;
  wire \$820 ;
  wire \$822 ;
  wire \$824 ;
  wire \$826 ;
  wire \$828 ;
  wire \$83 ;
  wire \$830 ;
  wire \$832 ;
  wire \$834 ;
  wire \$836 ;
  wire \$838 ;
  wire \$840 ;
  wire \$842 ;
  wire \$844 ;
  wire \$846 ;
  wire \$848 ;
  wire \$85 ;
  wire \$850 ;
  wire \$852 ;
  wire \$854 ;
  wire \$856 ;
  wire \$858 ;
  wire \$860 ;
  wire \$862 ;
  wire \$864 ;
  wire \$866 ;
  wire \$868 ;
  wire \$87 ;
  wire \$870 ;
  wire \$872 ;
  wire \$874 ;
  wire \$876 ;
  wire \$878 ;
  wire \$880 ;
  wire \$882 ;
  wire \$884 ;
  wire \$886 ;
  wire \$888 ;
  wire \$89 ;
  wire \$890 ;
  wire \$892 ;
  wire \$894 ;
  wire \$896 ;
  wire \$898 ;
  wire \$900 ;
  wire \$902 ;
  wire \$904 ;
  wire \$906 ;
  wire \$908 ;
  wire \$91 ;
  wire \$910 ;
  wire \$912 ;
  wire \$914 ;
  wire \$916 ;
  wire \$918 ;
  wire \$920 ;
  wire \$922 ;
  wire [34:0] \$924 ;
  wire [32:0] \$925 ;
  wire [33:0] \$927 ;
  wire [34:0] \$929 ;
  wire \$93 ;
  wire \$931 ;
  wire \$933 ;
  wire \$935 ;
  wire \$937 ;
  wire \$939 ;
  wire \$941 ;
  wire \$943 ;
  wire \$945 ;
  wire \$947 ;
  wire \$949 ;
  wire \$95 ;
  wire \$951 ;
  wire \$953 ;
  wire \$955 ;
  wire \$957 ;
  wire \$959 ;
  wire \$961 ;
  wire \$963 ;
  wire \$965 ;
  wire \$967 ;
  wire \$969 ;
  wire \$97 ;
  wire \$971 ;
  wire \$973 ;
  wire \$975 ;
  wire \$977 ;
  wire \$979 ;
  wire \$981 ;
  wire \$983 ;
  wire \$985 ;
  wire [2:0] \$987 ;
  wire [2:0] \$988 ;
  wire \$99 ;
  wire \$990 ;
  wire \$992 ;
  wire \$994 ;
  wire \$996 ;
  wire \$998 ;
  reg [31:0] bigK;
  reg [31:0] bp_a = 32'd0;
  reg [31:0] \bp_a$next ;
  reg [31:0] bp_b = 32'd0;
  reg [31:0] \bp_b$next ;
  reg [31:0] bp_c = 32'd0;
  reg [31:0] \bp_c$next ;
  reg [31:0] bp_d = 32'd0;
  reg [31:0] \bp_d$next ;
  reg [31:0] bp_e = 32'd0;
  reg [31:0] \bp_e$next ;
  reg [31:0] bp_f = 32'd0;
  reg [31:0] \bp_f$next ;
  reg [31:0] bp_g = 32'd0;
  reg [31:0] \bp_g$next ;
  reg [31:0] bp_h = 32'd0;
  reg [31:0] \bp_h$next ;
  reg bp_outrdy = 1'h0;
  reg \bp_outrdy$next ;
  (* enum_base_type = "BlockProcessorState" *)
  (* enum_value_0000 = "PowerUp" *)
  (* enum_value_0001 = "NewMessageBegin" *)
  (* enum_value_0010 = "NewBlockBegin" *)
  (* enum_value_0011 = "WaitForReady" *)
  (* enum_value_0100 = "ValueSnapShot" *)
  (* enum_value_0101 = "ProcessBlockUnit" *)
  (* enum_value_0110 = "CheckBlockDone" *)
  (* enum_value_0111 = "ProcessBlockDone" *)
  (* enum_value_1000 = "HashReady" *)
  reg [3:0] bp_procst = 4'h0;
  reg [3:0] \bp_procst$next ;
  output busy;
  reg busy = 1'h0;
  reg \busy$next ;
  wire [31:0] ch_ch_out;
  wire [31:0] ch_ch_x;
  wire [31:0] ch_ch_y;
  wire [31:0] ch_ch_z;
  reg checkedResults = 1'h0;
  reg \checkedResults$next ;
  input clk;
  wire clk;
  reg [31:0] currentResult = 32'd0;
  reg [31:0] \currentResult$next ;
  reg [31:0] debug_sig = 32'd0;
  reg [31:0] \debug_sig$next ;
  reg [3:0] delayCount = 4'h0;
  reg [3:0] \delayCount$next ;
  reg doProcessBlock = 1'h0;
  reg \doProcessBlock$next ;
  reg [31:0] hbuf0 = 32'd0;
  reg [31:0] \hbuf0$next ;
  reg [31:0] hbuf1 = 32'd0;
  reg [31:0] \hbuf1$next ;
  reg [31:0] hbuf2 = 32'd0;
  reg [31:0] \hbuf2$next ;
  reg [31:0] hbuf3 = 32'd0;
  reg [31:0] \hbuf3$next ;
  reg [31:0] hbuf4 = 32'd0;
  reg [31:0] \hbuf4$next ;
  reg [31:0] hbuf5 = 32'd0;
  reg [31:0] \hbuf5$next ;
  reg [31:0] hbuf6 = 32'd0;
  reg [31:0] \hbuf6$next ;
  reg [31:0] hbuf7 = 32'd0;
  reg [31:0] \hbuf7$next ;
  reg [511:0] hist = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  reg [511:0] \hist$next ;
  reg [3:0] in0 = 4'h0;
  reg [3:0] \in0$next ;
  reg [3:0] in1 = 4'h0;
  reg [3:0] \in1$next ;
  reg [3:0] in2 = 4'h0;
  reg [3:0] \in2$next ;
  reg [3:0] in3 = 4'h0;
  reg [3:0] \in3$next ;
  reg [3:0] in4 = 4'h0;
  reg [3:0] \in4$next ;
  reg [3:0] in5 = 4'h0;
  reg [3:0] \in5$next ;
  reg [3:0] in6 = 4'h0;
  reg [3:0] \in6$next ;
  reg [3:0] in7 = 4'h0;
  reg [3:0] \in7$next ;
  input [3:0] inNibble;
  wire [3:0] inNibble;
  wire [31:0] inWord;
  input inputReady;
  wire inputReady;
  reg inputSeen = 1'h0;
  reg \inputSeen$next ;
  reg [6:0] lastCount = 7'h00;
  reg [6:0] \lastCount$next ;
  reg [31:0] lastResult = 32'd0;
  reg [31:0] \lastResult$next ;
  reg [31:0] lastVal = 32'd0;
  reg [31:0] \lastVal$next ;
  reg myOutReady;
  reg newMessage = 1'h0;
  reg \newMessage$next ;
  reg [7:0] nibbleCount = 8'h00;
  reg [7:0] \nibbleCount$next ;
  reg [3:0] nibbleShift = 4'h0;
  reg [3:0] \nibbleShift$next ;
  output [3:0] nres_out;
  reg [3:0] nres_out = 4'h0;
  reg [3:0] \nres_out$next ;
  reg [31:0] opT1Output = 32'd0;
  reg [31:0] \opT1Output$next ;
  reg [31:0] opT2Output = 32'd0;
  reg [31:0] \opT2Output$next ;
  wire result;
  reg [5:0] resultOutputNibble = 6'h00;
  reg [5:0] \resultOutputNibble$next ;
  wire [31:0] rot1_rot1_out;
  wire [31:0] rot1_rot1_x;
  input rst;
  wire rst;
  wire [31:0] s0_s0_out;
  wire [31:0] s0_s0_x;
  wire [31:0] s1_s1_out;
  wire [31:0] s1_s1_x;
  reg [31:0] \sbuf-1  = 32'd0;
  reg [31:0] \sbuf-1$next ;
  reg [31:0] \sbuf-10  = 32'd0;
  reg [31:0] \sbuf-10$next ;
  reg [31:0] \sbuf-11  = 32'd0;
  reg [31:0] \sbuf-11$next ;
  reg [31:0] \sbuf-12  = 32'd0;
  reg [31:0] \sbuf-12$next ;
  reg [31:0] \sbuf-13  = 32'd0;
  reg [31:0] \sbuf-13$next ;
  reg [31:0] \sbuf-14  = 32'd0;
  reg [31:0] \sbuf-14$next ;
  reg [31:0] \sbuf-15  = 32'd0;
  reg [31:0] \sbuf-15$next ;
  reg [31:0] \sbuf-2  = 32'd0;
  reg [31:0] \sbuf-2$next ;
  reg [31:0] \sbuf-3  = 32'd0;
  reg [31:0] \sbuf-3$next ;
  reg [31:0] \sbuf-4  = 32'd0;
  reg [31:0] \sbuf-4$next ;
  reg [31:0] \sbuf-5  = 32'd0;
  reg [31:0] \sbuf-5$next ;
  reg [31:0] \sbuf-6  = 32'd0;
  reg [31:0] \sbuf-6$next ;
  reg [31:0] \sbuf-7  = 32'd0;
  reg [31:0] \sbuf-7$next ;
  reg [31:0] \sbuf-8  = 32'd0;
  reg [31:0] \sbuf-8$next ;
  reg [31:0] \sbuf-9  = 32'd0;
  reg [31:0] \sbuf-9$next ;
  reg [8:0] shiftCount = 9'h000;
  reg [8:0] \shiftCount$next ;
  reg [6:0] t1_count = 7'h00;
  reg [6:0] \t1_count$next ;
  wire [31:0] t1_e;
  wire [31:0] t1_f;
  wire [31:0] t1_g;
  wire [31:0] t1_h;
  wire [31:0] t1_out;
  wire t1_outrdy;
  wire [31:0] t2_t2_a;
  wire [31:0] t2_t2_b;
  wire [31:0] t2_t2_c;
  wire [31:0] t2_t2_out;
  reg thisIsLastUnitInBlock = 1'h0;
  reg \thisIsLastUnitInBlock$next ;
  reg [1:0] tickDelay = 2'h0;
  reg [1:0] \tickDelay$next ;
  reg [4:0] wordCount = 5'h00;
  reg [4:0] \wordCount$next ;
  wire [5:0] wt_count;
  reg [5:0] wt_lastcnt = 6'h00;
  reg [5:0] \wt_lastcnt$next ;
  reg [31:0] wt_out = 32'd0;
  reg [31:0] \wt_out$next ;
  reg wt_outrdy = 1'h0;
  reg \wt_outrdy$next ;
  wire [31:0] wt_res;
  assign \$99  = resultOutputNibble == 6'h20;
  assign \$1000  = wt_count < 5'h10;
  assign \$1002  = wt_count > wt_lastcnt;
  assign \$1004  = ! tickDelay;
  assign \$1006  = wt_count > 5'h10;
  assign \$1009  = shiftCount + 1'h1;
  assign \$1011  = wt_count < 5'h10;
  assign \$1013  = wt_count > wt_lastcnt;
  assign \$1015  = ! tickDelay;
  assign \$1017  = wt_count > 5'h10;
  assign \$101  = resultOutputNibble == 6'h21;
  assign \$1019  = wt_count < 5'h10;
  assign \$1021  = wt_count > wt_lastcnt;
  assign \$1023  = ! tickDelay;
  assign \$1025  = wt_count > 5'h10;
  assign \$1027  = wt_count < 5'h10;
  assign \$1029  = wt_count > wt_lastcnt;
  assign \$1031  = ! tickDelay;
  assign \$1033  = wt_count > 5'h10;
  assign \$1035  = wt_count < 5'h10;
  assign \$1037  = wt_count > wt_lastcnt;
  assign \$103  = resultOutputNibble == 6'h22;
  assign \$1039  = ! tickDelay;
  assign \$1041  = wt_count > 5'h10;
  assign \$1043  = wt_count < 5'h10;
  assign \$1045  = wt_count > wt_lastcnt;
  assign \$1047  = ! tickDelay;
  assign \$1049  = wt_count > 5'h10;
  assign \$1051  = wt_count < 5'h10;
  assign \$1053  = wt_count > wt_lastcnt;
  assign \$1055  = ! tickDelay;
  assign \$1057  = wt_count > 5'h10;
  assign \$105  = resultOutputNibble == 6'h23;
  assign \$1059  = wt_count < 5'h10;
  assign \$1061  = wt_count > wt_lastcnt;
  assign \$1063  = ! tickDelay;
  assign \$1065  = wt_count > 5'h10;
  assign \$1067  = wt_count < 5'h10;
  assign \$1069  = wt_count > wt_lastcnt;
  assign \$1071  = ! tickDelay;
  assign \$1073  = wt_count > 5'h10;
  assign \$1075  = wt_count < 5'h10;
  assign \$1077  = wt_count > wt_lastcnt;
  assign \$107  = resultOutputNibble == 6'h24;
  assign \$1079  = ! tickDelay;
  assign \$1081  = wt_count > 5'h10;
  assign \$1083  = wt_count < 5'h10;
  assign \$1085  = wt_count > wt_lastcnt;
  assign \$1087  = ! tickDelay;
  assign \$1089  = wt_count > 5'h10;
  assign \$1091  = wt_count < 5'h10;
  assign \$1093  = wt_count > wt_lastcnt;
  assign \$1095  = ! tickDelay;
  assign \$1097  = wt_count > 5'h10;
  assign \$10  = \$6  | \$8 ;
  assign \$109  = resultOutputNibble == 6'h25;
  assign \$1099  = wt_count < 5'h10;
  assign \$1101  = wt_count > wt_lastcnt;
  assign \$1103  = ! tickDelay;
  assign \$1105  = wt_count > 5'h10;
  assign \$1107  = wt_count < 5'h10;
  assign \$1109  = wt_count > wt_lastcnt;
  assign \$1111  = ! tickDelay;
  assign \$1113  = wt_count > 5'h10;
  assign \$1115  = wt_count < 5'h10;
  assign \$1117  = wt_count > wt_lastcnt;
  assign \$111  = resultOutputNibble == 6'h26;
  assign \$1119  = ! tickDelay;
  assign \$1121  = wt_count > 5'h10;
  assign \$1123  = wt_count < 5'h10;
  assign \$1125  = wt_count > wt_lastcnt;
  assign \$1127  = ! tickDelay;
  assign \$1129  = wt_count > 5'h10;
  assign \$1131  = wt_count < 5'h10;
  assign \$1133  = wt_count > wt_lastcnt;
  assign \$1135  = ! tickDelay;
  assign \$1137  = wt_count > 5'h10;
  assign \$113  = resultOutputNibble == 6'h27;
  assign \$1140  = debug_sig + 1'h1;
  assign \$1142  = wt_count < 5'h10;
  assign \$1144  = wt_count > wt_lastcnt;
  assign \$1146  = tickDelay == 1'h1;
  assign \$1148  = wt_count < 5'h10;
  assign \$1150  = wt_count > wt_lastcnt;
  assign \$1152  = tickDelay == 1'h1;
  always @(posedge clk)
    resultOutputNibble <= \resultOutputNibble$next ;
  always @(posedge clk)
    doProcessBlock <= \doProcessBlock$next ;
  always @(posedge clk)
    busy <= \busy$next ;
  always @(posedge clk)
    checkedResults <= \checkedResults$next ;
  always @(posedge clk)
    nres_out <= \nres_out$next ;
  always @(posedge clk)
    newMessage <= \newMessage$next ;
  assign \$115  = resultOutputNibble == 6'h28;
  always @(posedge clk)
    in0 <= \in0$next ;
  always @(posedge clk)
    in1 <= \in1$next ;
  always @(posedge clk)
    in2 <= \in2$next ;
  always @(posedge clk)
    in3 <= \in3$next ;
  always @(posedge clk)
    in4 <= \in4$next ;
  always @(posedge clk)
    in5 <= \in5$next ;
  always @(posedge clk)
    in6 <= \in6$next ;
  always @(posedge clk)
    in7 <= \in7$next ;
  always @(posedge clk)
    inputSeen <= \inputSeen$next ;
  always @(posedge clk)
    nibbleShift <= \nibbleShift$next ;
  always @(posedge clk)
    nibbleCount <= \nibbleCount$next ;
  always @(posedge clk)
    hist <= \hist$next ;
  always @(posedge clk)
    wordCount <= \wordCount$next ;
  always @(posedge clk)
    bp_procst <= \bp_procst$next ;
  always @(posedge clk)
    t1_count <= \t1_count$next ;
  always @(posedge clk)
    hbuf0 <= \hbuf0$next ;
  always @(posedge clk)
    hbuf1 <= \hbuf1$next ;
  always @(posedge clk)
    hbuf2 <= \hbuf2$next ;
  always @(posedge clk)
    hbuf3 <= \hbuf3$next ;
  always @(posedge clk)
    hbuf4 <= \hbuf4$next ;
  assign \$117  = resultOutputNibble == 6'h29;
  always @(posedge clk)
    hbuf5 <= \hbuf5$next ;
  always @(posedge clk)
    hbuf6 <= \hbuf6$next ;
  always @(posedge clk)
    hbuf7 <= \hbuf7$next ;
  always @(posedge clk)
    thisIsLastUnitInBlock <= \thisIsLastUnitInBlock$next ;
  always @(posedge clk)
    bp_outrdy <= \bp_outrdy$next ;
  always @(posedge clk)
    bp_a <= \bp_a$next ;
  always @(posedge clk)
    bp_b <= \bp_b$next ;
  always @(posedge clk)
    bp_c <= \bp_c$next ;
  always @(posedge clk)
    bp_d <= \bp_d$next ;
  always @(posedge clk)
    bp_e <= \bp_e$next ;
  always @(posedge clk)
    bp_f <= \bp_f$next ;
  always @(posedge clk)
    bp_g <= \bp_g$next ;
  always @(posedge clk)
    bp_h <= \bp_h$next ;
  always @(posedge clk)
    opT1Output <= \opT1Output$next ;
  always @(posedge clk)
    opT2Output <= \opT2Output$next ;
  always @(posedge clk)
    delayCount <= \delayCount$next ;
  always @(posedge clk)
    lastCount <= \lastCount$next ;
  always @(posedge clk)
    wt_lastcnt <= \wt_lastcnt$next ;
  always @(posedge clk)
    wt_outrdy <= \wt_outrdy$next ;
  always @(posedge clk)
    wt_out <= \wt_out$next ;
  assign \$119  = resultOutputNibble == 6'h2a;
  always @(posedge clk)
    tickDelay <= \tickDelay$next ;
  always @(posedge clk)
    lastVal <= \lastVal$next ;
  always @(posedge clk)
    shiftCount <= \shiftCount$next ;
  always @(posedge clk)
    \sbuf-1  <= \sbuf-1$next ;
  always @(posedge clk)
    \sbuf-2  <= \sbuf-2$next ;
  always @(posedge clk)
    \sbuf-3  <= \sbuf-3$next ;
  always @(posedge clk)
    \sbuf-4  <= \sbuf-4$next ;
  always @(posedge clk)
    \sbuf-5  <= \sbuf-5$next ;
  always @(posedge clk)
    \sbuf-6  <= \sbuf-6$next ;
  always @(posedge clk)
    \sbuf-7  <= \sbuf-7$next ;
  always @(posedge clk)
    \sbuf-8  <= \sbuf-8$next ;
  always @(posedge clk)
    \sbuf-9  <= \sbuf-9$next ;
  always @(posedge clk)
    \sbuf-10  <= \sbuf-10$next ;
  always @(posedge clk)
    \sbuf-11  <= \sbuf-11$next ;
  always @(posedge clk)
    \sbuf-12  <= \sbuf-12$next ;
  always @(posedge clk)
    \sbuf-13  <= \sbuf-13$next ;
  always @(posedge clk)
    \sbuf-14  <= \sbuf-14$next ;
  always @(posedge clk)
    \sbuf-15  <= \sbuf-15$next ;
  always @(posedge clk)
    debug_sig <= \debug_sig$next ;
  always @(posedge clk)
    lastResult <= \lastResult$next ;
  assign \$121  = resultOutputNibble == 6'h2b;
  always @(posedge clk)
    currentResult <= \currentResult$next ;
  assign \$123  = resultOutputNibble == 6'h2c;
  assign \$125  = resultOutputNibble == 6'h2d;
  assign \$127  = resultOutputNibble == 6'h2e;
  assign \$129  = resultOutputNibble == 6'h2f;
  assign \$131  = resultOutputNibble == 6'h30;
  assign \$133  = resultOutputNibble == 6'h31;
  assign \$135  = resultOutputNibble == 6'h32;
  assign \$137  = resultOutputNibble == 6'h33;
  assign \$139  = resultOutputNibble == 6'h34;
  assign \$141  = resultOutputNibble == 6'h35;
  assign \$143  = resultOutputNibble == 6'h36;
  assign \$145  = resultOutputNibble == 6'h37;
  assign \$147  = resultOutputNibble == 6'h38;
  assign \$14  = \$10  | \$12 ;
  assign \$149  = resultOutputNibble == 6'h39;
  assign \$151  = resultOutputNibble == 6'h3a;
  assign \$153  = resultOutputNibble == 6'h3b;
  assign \$155  = resultOutputNibble == 6'h3c;
  assign \$157  = resultOutputNibble == 6'h3d;
  assign \$159  = resultOutputNibble == 6'h3e;
  assign \$161  = resultOutputNibble == 6'h3f;
  assign \$163  = nibbleCount < 8'h80;
  assign \$165  = ! resultOutputNibble;
  assign \$168  = hbuf0 & 32'd4026531840;
  assign \$172  = resultOutputNibble == 1'h1;
  assign \$175  = hbuf0 & 28'hf000000;
  assign \$179  = resultOutputNibble == 2'h2;
  assign \$182  = hbuf0 & 24'hf00000;
  assign \$186  = resultOutputNibble == 2'h3;
  assign \$18  = \$14  | \$16 ;
  assign \$189  = hbuf0 & 20'hf0000;
  assign \$193  = resultOutputNibble == 3'h4;
  assign \$196  = hbuf0 & 16'hf000;
  assign \$200  = resultOutputNibble == 3'h5;
  assign \$203  = hbuf0 & 12'hf00;
  assign \$207  = resultOutputNibble == 3'h6;
  assign \$210  = hbuf0 & 8'hf0;
  assign \$214  = resultOutputNibble == 3'h7;
  assign \$217  = hbuf0 & 4'hf;
  assign \$221  = resultOutputNibble == 4'h8;
  assign \$224  = hbuf1 & 32'd4026531840;
  assign \$228  = resultOutputNibble == 4'h9;
  assign \$22  = \$18  | \$20 ;
  assign \$231  = hbuf1 & 28'hf000000;
  assign \$235  = resultOutputNibble == 4'ha;
  assign \$238  = hbuf1 & 24'hf00000;
  assign \$242  = resultOutputNibble == 4'hb;
  assign \$245  = hbuf1 & 20'hf0000;
  assign \$249  = resultOutputNibble == 4'hc;
  assign \$252  = hbuf1 & 16'hf000;
  assign \$256  = resultOutputNibble == 4'hd;
  assign \$259  = hbuf1 & 12'hf00;
  assign \$263  = resultOutputNibble == 4'he;
  assign \$266  = hbuf1 & 8'hf0;
  assign \$26  = \$22  | \$24 ;
  assign \$270  = resultOutputNibble == 4'hf;
  assign \$273  = hbuf1 & 4'hf;
  assign \$277  = resultOutputNibble == 5'h10;
  assign \$280  = hbuf2 & 32'd4026531840;
  assign \$284  = resultOutputNibble == 5'h11;
  assign \$287  = hbuf2 & 28'hf000000;
  assign \$28  = \$26  | in7;
  assign \$291  = resultOutputNibble == 5'h12;
  assign \$294  = hbuf2 & 24'hf00000;
  assign \$298  = resultOutputNibble == 5'h13;
  assign \$301  = hbuf2 & 20'hf0000;
  assign \$305  = resultOutputNibble == 5'h14;
  assign \$308  = hbuf2 & 16'hf000;
  assign \$312  = resultOutputNibble == 5'h15;
  assign \$315  = hbuf2 & 12'hf00;
  assign \$31  = resultOutputNibble + 1'h1;
  assign \$319  = resultOutputNibble == 5'h16;
  assign \$322  = hbuf2 & 8'hf0;
  assign \$326  = resultOutputNibble == 5'h17;
  assign \$329  = hbuf2 & 4'hf;
  assign \$333  = resultOutputNibble == 5'h18;
  assign \$336  = hbuf3 & 32'd4026531840;
  assign \$33  = nibbleCount < 8'h80;
  assign \$340  = resultOutputNibble == 5'h19;
  assign \$343  = hbuf3 & 28'hf000000;
  assign \$347  = resultOutputNibble == 5'h1a;
  assign \$350  = hbuf3 & 24'hf00000;
  assign \$354  = resultOutputNibble == 5'h1b;
  assign \$357  = hbuf3 & 20'hf0000;
  assign \$35  = ! resultOutputNibble;
  assign \$361  = resultOutputNibble == 5'h1c;
  assign \$364  = hbuf3 & 16'hf000;
  assign \$368  = resultOutputNibble == 5'h1d;
  assign \$371  = hbuf3 & 12'hf00;
  assign \$375  = resultOutputNibble == 5'h1e;
  assign \$378  = hbuf3 & 8'hf0;
  assign \$37  = resultOutputNibble == 1'h1;
  assign \$382  = resultOutputNibble == 5'h1f;
  assign \$385  = hbuf3 & 4'hf;
  assign \$389  = resultOutputNibble == 6'h20;
  assign \$392  = hbuf4 & 32'd4026531840;
  assign \$396  = resultOutputNibble == 6'h21;
  assign \$39  = resultOutputNibble == 2'h2;
  assign \$399  = hbuf4 & 28'hf000000;
  assign \$403  = resultOutputNibble == 6'h22;
  assign \$406  = hbuf4 & 24'hf00000;
  assign \$410  = resultOutputNibble == 6'h23;
  assign \$413  = hbuf4 & 20'hf0000;
  assign \$417  = resultOutputNibble == 6'h24;
  assign \$41  = resultOutputNibble == 2'h3;
  assign \$420  = hbuf4 & 16'hf000;
  assign \$424  = resultOutputNibble == 6'h25;
  assign \$427  = hbuf4 & 12'hf00;
  assign \$431  = resultOutputNibble == 6'h26;
  assign \$434  = hbuf4 & 8'hf0;
  assign \$438  = resultOutputNibble == 6'h27;
  assign \$43  = resultOutputNibble == 3'h4;
  assign \$441  = hbuf4 & 4'hf;
  assign \$445  = resultOutputNibble == 6'h28;
  assign \$448  = hbuf5 & 32'd4026531840;
  assign \$452  = resultOutputNibble == 6'h29;
  assign \$455  = hbuf5 & 28'hf000000;
  assign \$45  = resultOutputNibble == 3'h5;
  assign \$459  = resultOutputNibble == 6'h2a;
  assign \$462  = hbuf5 & 24'hf00000;
  assign \$466  = resultOutputNibble == 6'h2b;
  assign \$469  = hbuf5 & 20'hf0000;
  assign \$473  = resultOutputNibble == 6'h2c;
  assign \$476  = hbuf5 & 16'hf000;
  assign \$47  = resultOutputNibble == 3'h6;
  assign \$480  = resultOutputNibble == 6'h2d;
  assign \$483  = hbuf5 & 12'hf00;
  assign \$487  = resultOutputNibble == 6'h2e;
  assign \$490  = hbuf5 & 8'hf0;
  assign \$494  = resultOutputNibble == 6'h2f;
  assign \$497  = hbuf5 & 4'hf;
  assign \$49  = resultOutputNibble == 3'h7;
  assign \$501  = resultOutputNibble == 6'h30;
  assign \$504  = hbuf6 & 32'd4026531840;
  assign \$508  = resultOutputNibble == 6'h31;
  assign \$511  = hbuf6 & 28'hf000000;
  assign \$515  = resultOutputNibble == 6'h32;
  assign \$518  = hbuf6 & 24'hf00000;
  assign \$51  = resultOutputNibble == 4'h8;
  assign \$522  = resultOutputNibble == 6'h33;
  assign \$525  = hbuf6 & 20'hf0000;
  assign \$529  = resultOutputNibble == 6'h34;
  assign \$532  = hbuf6 & 16'hf000;
  assign \$536  = resultOutputNibble == 6'h35;
  assign \$53  = resultOutputNibble == 4'h9;
  assign \$539  = hbuf6 & 12'hf00;
  assign \$543  = resultOutputNibble == 6'h36;
  assign \$546  = hbuf6 & 8'hf0;
  assign \$550  = resultOutputNibble == 6'h37;
  assign \$553  = hbuf6 & 4'hf;
  assign \$557  = resultOutputNibble == 6'h38;
  assign \$55  = resultOutputNibble == 4'ha;
  assign \$560  = hbuf7 & 32'd4026531840;
  assign \$564  = resultOutputNibble == 6'h39;
  assign \$567  = hbuf7 & 28'hf000000;
  assign \$571  = resultOutputNibble == 6'h3a;
  assign \$574  = hbuf7 & 24'hf00000;
  assign \$578  = resultOutputNibble == 6'h3b;
  assign \$57  = resultOutputNibble == 4'hb;
  assign \$581  = hbuf7 & 20'hf0000;
  assign \$585  = resultOutputNibble == 6'h3c;
  assign \$588  = hbuf7 & 16'hf000;
  assign \$592  = resultOutputNibble == 6'h3d;
  assign \$595  = hbuf7 & 12'hf00;
  assign \$59  = resultOutputNibble == 4'hc;
  assign \$599  = resultOutputNibble == 6'h3e;
  assign \$602  = hbuf7 & 8'hf0;
  assign \$606  = resultOutputNibble == 6'h3f;
  assign \$609  = hbuf7 & 4'hf;
  assign \$613  = nibbleCount < 8'h80;
  assign \$615  = ~ inputSeen;
  assign \$617  = ! nibbleShift;
  assign \$61  = resultOutputNibble == 4'hd;
  assign \$619  = nibbleCount < 8'h80;
  assign \$621  = ~ inputSeen;
  assign \$623  = nibbleShift == 1'h1;
  assign \$625  = nibbleCount < 8'h80;
  assign \$627  = ~ inputSeen;
  assign \$629  = nibbleShift == 2'h2;
  assign \$631  = nibbleCount < 8'h80;
  assign \$633  = ~ inputSeen;
  assign \$635  = nibbleShift == 2'h3;
  assign \$637  = nibbleCount < 8'h80;
  assign \$63  = resultOutputNibble == 4'he;
  assign \$639  = ~ inputSeen;
  assign \$641  = nibbleShift == 3'h4;
  assign \$643  = nibbleCount < 8'h80;
  assign \$645  = ~ inputSeen;
  assign \$647  = nibbleShift == 3'h5;
  assign \$649  = nibbleCount < 8'h80;
  assign \$651  = ~ inputSeen;
  assign \$653  = nibbleShift == 3'h6;
  assign \$655  = nibbleCount < 8'h80;
  assign \$657  = ~ inputSeen;
  assign \$65  = resultOutputNibble == 4'hf;
  assign \$659  = nibbleShift == 3'h7;
  assign \$661  = nibbleCount < 8'h80;
  assign \$663  = ~ inputSeen;
  assign \$665  = nibbleCount < 8'h80;
  assign \$667  = ~ inputSeen;
  assign \$670  = nibbleShift + 1'h1;
  assign \$672  = nibbleShift == 4'h8;
  assign \$674  = nibbleCount < 8'h80;
  assign \$676  = ~ inputSeen;
  assign \$67  = resultOutputNibble == 5'h10;
  assign \$679  = nibbleCount + 1'h1;
  assign \$681  = nibbleCount < 8'h80;
  assign \$683  = nibbleShift == 4'h8;
  assign \$685  = ! wordCount;
  assign \$687  = wordCount == 1'h1;
  assign \$689  = wordCount == 2'h2;
  assign \$691  = wordCount == 2'h3;
  assign \$693  = wordCount == 3'h4;
  assign \$695  = wordCount == 3'h5;
  assign \$697  = wordCount == 3'h6;
  assign \$6  = \$2  | \$4 ;
  assign \$69  = resultOutputNibble == 5'h11;
  assign \$699  = wordCount == 3'h7;
  assign \$701  = wordCount == 4'h8;
  assign \$703  = wordCount == 4'h9;
  assign \$705  = wordCount == 4'ha;
  assign \$707  = wordCount == 4'hb;
  assign \$709  = wordCount == 4'hc;
  assign \$711  = wordCount == 4'hd;
  assign \$713  = wordCount == 4'he;
  assign \$715  = wordCount == 4'hf;
  assign \$717  = wt_count < 5'h10;
  assign \$71  = resultOutputNibble == 5'h12;
  assign \$719  = wt_count > wt_lastcnt;
  assign \$721  = ! tickDelay;
  assign \$723  = wt_count > 5'h10;
  assign \$728  = \$726  | currentResult;
  assign \$730  = nibbleCount < 8'h80;
  assign \$732  = nibbleShift == 4'h8;
  assign \$735  = wordCount + 1'h1;
  assign \$737  = ~ doProcessBlock;
  assign \$73  = resultOutputNibble == 5'h13;
  assign \$740  = t1_count + 1'h1;
  assign \$743  = hbuf0 + bp_a;
  assign \$746  = hbuf1 + bp_b;
  assign \$749  = hbuf2 + bp_c;
  assign \$752  = hbuf3 + bp_d;
  assign \$755  = hbuf4 + bp_e;
  assign \$758  = hbuf5 + bp_f;
  assign \$75  = resultOutputNibble == 5'h14;
  assign \$761  = hbuf6 + bp_g;
  assign \$764  = hbuf7 + bp_h;
  assign \$766  = t1_count == 6'h3f;
  assign \$768  = ~ doProcessBlock;
  assign \$771  = opT1Output + opT2Output;
  assign \$774  = bp_d + opT1Output;
  assign \$776  = lastCount != t1_count;
  assign \$778  = delayCount < 3'h4;
  assign \$77  = resultOutputNibble == 5'h15;
  assign \$781  = delayCount + 1'h1;
  assign \$783  = lastCount != t1_count;
  assign \$785  = delayCount < 3'h4;
  assign \$788  = t1_h + rot1_rot1_out;
  assign \$790  = \$788  + ch_ch_out;
  assign \$792  = \$790  + bigK;
  assign \$794  = \$792  + wt_out;
  assign \$796  = ! t1_count;
  assign \$798  = t1_count == 1'h1;
  assign \$79  = resultOutputNibble == 5'h16;
  assign \$800  = t1_count == 2'h2;
  assign \$802  = t1_count == 2'h3;
  assign \$804  = t1_count == 3'h4;
  assign \$806  = t1_count == 3'h5;
  assign \$808  = t1_count == 3'h6;
  assign \$810  = t1_count == 3'h7;
  assign \$812  = t1_count == 4'h8;
  assign \$814  = t1_count == 4'h9;
  assign \$816  = t1_count == 4'ha;
  assign \$818  = t1_count == 4'hb;
  assign \$81  = resultOutputNibble == 5'h17;
  assign \$820  = t1_count == 4'hc;
  assign \$822  = t1_count == 4'hd;
  assign \$824  = t1_count == 4'he;
  assign \$826  = t1_count == 4'hf;
  assign \$828  = t1_count == 5'h10;
  assign \$830  = t1_count == 5'h11;
  assign \$832  = t1_count == 5'h12;
  assign \$834  = t1_count == 5'h13;
  assign \$836  = t1_count == 5'h14;
  assign \$838  = t1_count == 5'h15;
  assign \$83  = resultOutputNibble == 5'h18;
  assign \$840  = t1_count == 5'h16;
  assign \$842  = t1_count == 5'h17;
  assign \$844  = t1_count == 5'h18;
  assign \$846  = t1_count == 5'h19;
  assign \$848  = t1_count == 5'h1a;
  assign \$850  = t1_count == 5'h1b;
  assign \$852  = t1_count == 5'h1c;
  assign \$854  = t1_count == 5'h1d;
  assign \$856  = t1_count == 5'h1e;
  assign \$858  = t1_count == 5'h1f;
  assign \$85  = resultOutputNibble == 5'h19;
  assign \$860  = t1_count == 6'h20;
  assign \$862  = t1_count == 6'h21;
  assign \$864  = t1_count == 6'h22;
  assign \$866  = t1_count == 6'h23;
  assign \$868  = t1_count == 6'h24;
  assign \$870  = t1_count == 6'h25;
  assign \$872  = t1_count == 6'h26;
  assign \$874  = t1_count == 6'h27;
  assign \$876  = t1_count == 6'h28;
  assign \$878  = t1_count == 6'h29;
  assign \$87  = resultOutputNibble == 5'h1a;
  assign \$880  = t1_count == 6'h2a;
  assign \$882  = t1_count == 6'h2b;
  assign \$884  = t1_count == 6'h2c;
  assign \$886  = t1_count == 6'h2d;
  assign \$888  = t1_count == 6'h2e;
  assign \$890  = t1_count == 6'h2f;
  assign \$892  = t1_count == 6'h30;
  assign \$894  = t1_count == 6'h31;
  assign \$896  = t1_count == 6'h32;
  assign \$898  = t1_count == 6'h33;
  assign \$89  = resultOutputNibble == 5'h1b;
  assign \$900  = t1_count == 6'h34;
  assign \$902  = t1_count == 6'h35;
  assign \$904  = t1_count == 6'h36;
  assign \$906  = t1_count == 6'h37;
  assign \$908  = t1_count == 6'h38;
  assign \$910  = t1_count == 6'h39;
  assign \$912  = t1_count == 6'h3a;
  assign \$914  = t1_count == 6'h3b;
  assign \$916  = t1_count == 6'h3c;
  assign \$918  = t1_count == 6'h3d;
  assign \$91  = resultOutputNibble == 5'h1c;
  assign \$920  = t1_count == 6'h3e;
  assign \$922  = t1_count == 6'h3f;
  assign \$925  = s1_s1_out + hist[223:192];
  assign \$927  = \$925  + s0_s0_out;
  assign \$929  = \$927  + hist[511:480];
  assign \$931  = wt_lastcnt > wt_count;
  assign \$933  = wt_count < 5'h10;
  assign \$935  = wt_count > wt_lastcnt;
  assign \$937  = tickDelay == 2'h2;
  assign \$93  = resultOutputNibble == 5'h1d;
  assign \$939  = wt_count < 5'h10;
  assign \$941  = wt_count > wt_lastcnt;
  assign \$943  = ! tickDelay;
  assign \$945  = tickDelay == 1'h1;
  assign \$947  = tickDelay == 2'h2;
  assign \$949  = wt_count < 5'h10;
  assign \$951  = ! wt_count;
  assign \$953  = wt_count == 1'h1;
  assign \$955  = wt_count == 2'h2;
  assign \$957  = wt_count == 2'h3;
  assign \$95  = resultOutputNibble == 5'h1e;
  assign \$959  = wt_count == 3'h4;
  assign \$961  = wt_count == 3'h5;
  assign \$963  = wt_count == 3'h6;
  assign \$965  = wt_count == 3'h7;
  assign \$967  = wt_count == 4'h8;
  assign \$969  = wt_count == 4'h9;
  assign \$971  = wt_count == 4'ha;
  assign \$973  = wt_count == 4'hb;
  assign \$975  = wt_count == 4'hc;
  assign \$977  = wt_count == 4'hd;
  assign \$97  = resultOutputNibble == 5'h1f;
  assign \$979  = wt_count == 4'he;
  assign \$981  = wt_count == 4'hf;
  assign \$983  = wt_count < 5'h10;
  assign \$985  = wt_count > wt_lastcnt;
  assign \$988  = tickDelay + 1'h1;
  assign \$990  = tickDelay == 2'h2;
  assign \$992  = wt_count < 5'h10;
  assign \$994  = wt_count > wt_lastcnt;
  assign \$996  = ! tickDelay;
  assign \$998  = wt_count > 5'h10;
  \buf  \buf  (
  );
  ch ch (
    .ch_out(ch_ch_out),
    .ch_x(ch_ch_x),
    .ch_y(ch_ch_y),
    .ch_z(ch_ch_z)
  );
  rot1 rot1 (
    .rot1_out(rot1_rot1_out),
    .rot1_x(rot1_rot1_x)
  );
  s0 s0 (
    .s0_out(s0_s0_out),
    .s0_x(s0_s0_x)
  );
  s1 s1 (
    .s1_out(s1_s1_out),
    .s1_x(s1_s1_x)
  );
  t2 t2 (
    .t2_a(t2_t2_a),
    .t2_b(t2_t2_b),
    .t2_c(t2_t2_c),
    .t2_out(t2_t2_out)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \resultOutputNibble$next  = resultOutputNibble;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          \resultOutputNibble$next  = \$31 [5:0];
      default:
          casez (checkedResults)
            1'h1:
                \resultOutputNibble$next  = 6'h00;
          endcase
    endcase
    casez (rst)
      1'h1:
          \resultOutputNibble$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in3$next  = in3;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$631 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$633 )
                        1'h1:
                            casez (\$635 )
                              1'h1:
                                  \in3$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in3$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in4$next  = in4;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$637 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$639 )
                        1'h1:
                            casez (\$641 )
                              1'h1:
                                  \in4$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in4$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in5$next  = in5;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$643 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$645 )
                        1'h1:
                            casez (\$647 )
                              1'h1:
                                  \in5$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in5$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in6$next  = in6;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$649 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$651 )
                        1'h1:
                            casez (\$653 )
                              1'h1:
                                  \in6$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in6$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in7$next  = in7;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$655 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$657 )
                        1'h1:
                            casez (\$659 )
                              1'h1:
                                  \in7$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in7$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \inputSeen$next  = inputSeen;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$661 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      casez (\$663 )
                        1'h1:
                            \inputSeen$next  = 1'h1;
                      endcase
                  default:
                      \inputSeen$next  = 1'h0;
                endcase
            default:
                casez (inputSeen)
                  1'h1:
                      \inputSeen$next  = 1'h0;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \inputSeen$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \nibbleShift$next  = nibbleShift;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$665 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      casez (\$667 )
                        1'h1:
                            \nibbleShift$next  = \$670 [3:0];
                      endcase
                  default:
                      casez (\$672 )
                        1'h1:
                            casez (inputSeen)
                              1'h1:
                                  \nibbleShift$next  = 4'h0;
                            endcase
                      endcase
                endcase
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      /* empty */;
                  default:
                      casez (bp_outrdy)
                        1'h1:
                            \nibbleShift$next  = 4'h0;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \nibbleShift$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \nibbleCount$next  = nibbleCount;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$674 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$676 )
                        1'h1:
                            \nibbleCount$next  = \$679 [7:0];
                      endcase
                endcase
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      /* empty */;
                  default:
                      casez (bp_outrdy)
                        1'h1:
                            \nibbleCount$next  = 8'h00;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \nibbleCount$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hist$next  = hist;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$681 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      /* empty */;
                  default:
                      casez (\$683 )
                        1'h1:
                            casez (inputSeen)
                              1'h1:
                                begin
                                  casez (\$685 )
                                    1'h1:
                                        \hist$next [511:480] = inWord;
                                  endcase
                                  casez (\$687 )
                                    1'h1:
                                        \hist$next [479:448] = inWord;
                                  endcase
                                  casez (\$689 )
                                    1'h1:
                                        \hist$next [447:416] = inWord;
                                  endcase
                                  casez (\$691 )
                                    1'h1:
                                        \hist$next [415:384] = inWord;
                                  endcase
                                  casez (\$693 )
                                    1'h1:
                                        \hist$next [383:352] = inWord;
                                  endcase
                                  casez (\$695 )
                                    1'h1:
                                        \hist$next [351:320] = inWord;
                                  endcase
                                  casez (\$697 )
                                    1'h1:
                                        \hist$next [319:288] = inWord;
                                  endcase
                                  casez (\$699 )
                                    1'h1:
                                        \hist$next [287:256] = inWord;
                                  endcase
                                  casez (\$701 )
                                    1'h1:
                                        \hist$next [255:224] = inWord;
                                  endcase
                                  casez (\$703 )
                                    1'h1:
                                        \hist$next [223:192] = inWord;
                                  endcase
                                  casez (\$705 )
                                    1'h1:
                                        \hist$next [191:160] = inWord;
                                  endcase
                                  casez (\$707 )
                                    1'h1:
                                        \hist$next [159:128] = inWord;
                                  endcase
                                  casez (\$709 )
                                    1'h1:
                                        \hist$next [127:96] = inWord;
                                  endcase
                                  casez (\$711 )
                                    1'h1:
                                        \hist$next [95:64] = inWord;
                                  endcase
                                  casez (\$713 )
                                    1'h1:
                                        \hist$next [63:32] = inWord;
                                  endcase
                                  casez (\$715 )
                                    1'h1:
                                        \hist$next [31:0] = inWord;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
            default:
                casez (inputSeen)
                  1'h1:
                      \hist$next [31:0] = inWord;
                endcase
          endcase
    endcase
    (* full_case = 32'd1 *)
    casez (\$717 )
      1'h1:
          /* empty */;
      default:
          casez (\$719 )
            1'h1:
                casez (\$721 )
                  1'h1:
                      casez (\$723 )
                        1'h1:
                            \hist$next  = \$728 [511:0];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \hist$next  = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \wordCount$next  = wordCount;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$730 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      /* empty */;
                  default:
                      casez (\$732 )
                        1'h1:
                            casez (inputSeen)
                              1'h1:
                                  \wordCount$next  = \$735 [4:0];
                            endcase
                      endcase
                endcase
            default:
                casez (inputSeen)
                  1'h1:
                      \wordCount$next  = 5'h00;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \wordCount$next  = 5'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \doProcessBlock$next  = doProcessBlock;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          \doProcessBlock$next  = 1'h0;
      default:
          (* full_case = 32'd1 *)
          casez (\$33 )
            1'h1:
                \doProcessBlock$next  = 1'h0;
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      /* empty */;
                  default:
                      \doProcessBlock$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \doProcessBlock$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_procst$next  = bp_procst;
    (* full_case = 32'd1 *)
    casez (bp_procst)
      4'h0:
          \bp_procst$next  = 4'h1;
      4'h1:
          \bp_procst$next  = 4'h2;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_procst$next  = 4'h3;
          endcase
      4'h3:
          casez (t1_outrdy)
            1'h1:
                \bp_procst$next  = 4'h4;
          endcase
      4'h4:
          \bp_procst$next  = 4'h5;
      4'h5:
          \bp_procst$next  = 4'h6;
      4'h6:
          (* full_case = 32'd1 *)
          casez (thisIsLastUnitInBlock)
            1'h1:
                \bp_procst$next  = 4'h7;
            default:
                \bp_procst$next  = 4'h3;
          endcase
      4'h7:
          \bp_procst$next  = 4'h8;
      4'h8:
          casez (\$737 )
            1'h1:
                \bp_procst$next  = 4'h2;
          endcase
      default:
          \bp_procst$next  = 4'h0;
    endcase
    casez (newMessage)
      1'h1:
          \bp_procst$next  = 4'h0;
    endcase
    casez (rst)
      1'h1:
          \bp_procst$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \t1_count$next  = t1_count;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \t1_count$next  = 7'h00;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \t1_count$next  = 7'h00;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \t1_count$next  = \$740 [6:0];
    endcase
    casez (rst)
      1'h1:
          \t1_count$next  = 7'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf0$next  = hbuf0;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf0$next  = 32'd1779033703;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf0$next  = \$743 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf0$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
        begin
          \busy$next  = 1'h1;
          casez (\$35 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$37 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$39 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$41 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$43 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$45 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$47 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$49 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$51 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$53 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$55 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$57 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$59 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$61 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$63 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$65 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$67 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$69 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$71 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$73 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$75 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$77 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$79 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$81 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$83 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$85 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$87 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$89 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$91 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$93 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$95 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$97 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$99 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$101 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$103 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$105 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$107 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$109 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$111 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$113 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$115 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$117 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$119 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$121 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$123 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$125 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$127 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$129 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$131 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$133 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$135 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$137 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$139 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$141 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$143 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$145 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$147 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$149 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$151 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$153 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$155 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$157 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$159 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
          casez (\$161 )
            1'h1:
                \busy$next  = 1'h0;
          endcase
        end
      default:
          (* full_case = 32'd1 *)
          casez (\$163 )
            1'h1:
                \busy$next  = 1'h0;
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      \busy$next  = 1'h1;
                  default:
                      (* full_case = 32'd1 *)
                      casez (bp_outrdy)
                        1'h1:
                            \busy$next  = 1'h0;
                        default:
                            \busy$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \busy$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf1$next  = hbuf1;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf1$next  = 32'd3144134277;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf1$next  = \$746 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf1$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf2$next  = hbuf2;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf2$next  = 32'd1013904242;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf2$next  = \$749 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf2$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf3$next  = hbuf3;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf3$next  = 32'd2773480762;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf3$next  = \$752 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf3$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf4$next  = hbuf4;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf4$next  = 32'd1359893119;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf4$next  = \$755 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf4$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf5$next  = hbuf5;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf5$next  = 32'd2600822924;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf5$next  = \$758 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf5$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf6$next  = hbuf6;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf6$next  = 32'd528734635;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf6$next  = \$761 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf6$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \hbuf7$next  = hbuf7;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          \hbuf7$next  = 32'd1541459225;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf7$next  = \$764 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf7$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \thisIsLastUnitInBlock$next  = thisIsLastUnitInBlock;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \thisIsLastUnitInBlock$next  = 1'h0;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          casez (\$766 )
            1'h1:
                \thisIsLastUnitInBlock$next  = 1'h1;
          endcase
    endcase
    casez (rst)
      1'h1:
          \thisIsLastUnitInBlock$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_outrdy$next  = bp_outrdy;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_outrdy$next  = 1'h0;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          /* empty */;
      4'h8:
        begin
          \bp_outrdy$next  = 1'h1;
          casez (\$768 )
            1'h1:
                \bp_outrdy$next  = 1'h0;
          endcase
        end
    endcase
    casez (rst)
      1'h1:
          \bp_outrdy$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_a$next  = bp_a;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_a$next  = hbuf0;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_a$next  = \$771 [31:0];
    endcase
    casez (rst)
      1'h1:
          \bp_a$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \checkedResults$next  = checkedResults;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          \checkedResults$next  = 1'h1;
      default:
          casez (checkedResults)
            1'h1:
                \checkedResults$next  = 1'h0;
          endcase
    endcase
    casez (rst)
      1'h1:
          \checkedResults$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_b$next  = bp_b;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_b$next  = hbuf1;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_b$next  = bp_a;
    endcase
    casez (rst)
      1'h1:
          \bp_b$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_c$next  = bp_c;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_c$next  = hbuf2;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_c$next  = bp_b;
    endcase
    casez (rst)
      1'h1:
          \bp_c$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_d$next  = bp_d;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_d$next  = hbuf3;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_d$next  = bp_c;
    endcase
    casez (rst)
      1'h1:
          \bp_d$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_e$next  = bp_e;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_e$next  = hbuf4;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_e$next  = \$774 [31:0];
    endcase
    casez (rst)
      1'h1:
          \bp_e$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_f$next  = bp_f;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_f$next  = hbuf5;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_f$next  = bp_e;
    endcase
    casez (rst)
      1'h1:
          \bp_f$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_g$next  = bp_g;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_g$next  = hbuf6;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_g$next  = bp_f;
    endcase
    casez (rst)
      1'h1:
          \bp_g$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \bp_h$next  = bp_h;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_h$next  = hbuf7;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_h$next  = bp_g;
    endcase
    casez (rst)
      1'h1:
          \bp_h$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \opT1Output$next  = opT1Output;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          \opT1Output$next  = t1_out;
    endcase
    casez (rst)
      1'h1:
          \opT1Output$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \opT2Output$next  = opT2Output;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          \opT2Output$next  = t2_t2_out;
    endcase
    casez (rst)
      1'h1:
          \opT2Output$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \delayCount$next  = delayCount;
    casez (\$776 )
      1'h1:
          \delayCount$next  = 4'h0;
    endcase
    casez (\$778 )
      1'h1:
          \delayCount$next  = \$781 [3:0];
    endcase
    casez (rst)
      1'h1:
          \delayCount$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \nres_out$next  = nres_out;
    casez (result)
      1'h1:
        begin
          casez (\$165 )
            1'h1:
                \nres_out$next  = \$170 [3:0];
          endcase
          casez (\$172 )
            1'h1:
                \nres_out$next  = \$177 [3:0];
          endcase
          casez (\$179 )
            1'h1:
                \nres_out$next  = \$184 [3:0];
          endcase
          casez (\$186 )
            1'h1:
                \nres_out$next  = \$191 [3:0];
          endcase
          casez (\$193 )
            1'h1:
                \nres_out$next  = \$198 [3:0];
          endcase
          casez (\$200 )
            1'h1:
                \nres_out$next  = \$205 [3:0];
          endcase
          casez (\$207 )
            1'h1:
                \nres_out$next  = \$212 [3:0];
          endcase
          casez (\$214 )
            1'h1:
                \nres_out$next  = \$219 [3:0];
          endcase
          casez (\$221 )
            1'h1:
                \nres_out$next  = \$226 [3:0];
          endcase
          casez (\$228 )
            1'h1:
                \nres_out$next  = \$233 [3:0];
          endcase
          casez (\$235 )
            1'h1:
                \nres_out$next  = \$240 [3:0];
          endcase
          casez (\$242 )
            1'h1:
                \nres_out$next  = \$247 [3:0];
          endcase
          casez (\$249 )
            1'h1:
                \nres_out$next  = \$254 [3:0];
          endcase
          casez (\$256 )
            1'h1:
                \nres_out$next  = \$261 [3:0];
          endcase
          casez (\$263 )
            1'h1:
                \nres_out$next  = \$268 [3:0];
          endcase
          casez (\$270 )
            1'h1:
                \nres_out$next  = \$275 [3:0];
          endcase
          casez (\$277 )
            1'h1:
                \nres_out$next  = \$282 [3:0];
          endcase
          casez (\$284 )
            1'h1:
                \nres_out$next  = \$289 [3:0];
          endcase
          casez (\$291 )
            1'h1:
                \nres_out$next  = \$296 [3:0];
          endcase
          casez (\$298 )
            1'h1:
                \nres_out$next  = \$303 [3:0];
          endcase
          casez (\$305 )
            1'h1:
                \nres_out$next  = \$310 [3:0];
          endcase
          casez (\$312 )
            1'h1:
                \nres_out$next  = \$317 [3:0];
          endcase
          casez (\$319 )
            1'h1:
                \nres_out$next  = \$324 [3:0];
          endcase
          casez (\$326 )
            1'h1:
                \nres_out$next  = \$331 [3:0];
          endcase
          casez (\$333 )
            1'h1:
                \nres_out$next  = \$338 [3:0];
          endcase
          casez (\$340 )
            1'h1:
                \nres_out$next  = \$345 [3:0];
          endcase
          casez (\$347 )
            1'h1:
                \nres_out$next  = \$352 [3:0];
          endcase
          casez (\$354 )
            1'h1:
                \nres_out$next  = \$359 [3:0];
          endcase
          casez (\$361 )
            1'h1:
                \nres_out$next  = \$366 [3:0];
          endcase
          casez (\$368 )
            1'h1:
                \nres_out$next  = \$373 [3:0];
          endcase
          casez (\$375 )
            1'h1:
                \nres_out$next  = \$380 [3:0];
          endcase
          casez (\$382 )
            1'h1:
                \nres_out$next  = \$387 [3:0];
          endcase
          casez (\$389 )
            1'h1:
                \nres_out$next  = \$394 [3:0];
          endcase
          casez (\$396 )
            1'h1:
                \nres_out$next  = \$401 [3:0];
          endcase
          casez (\$403 )
            1'h1:
                \nres_out$next  = \$408 [3:0];
          endcase
          casez (\$410 )
            1'h1:
                \nres_out$next  = \$415 [3:0];
          endcase
          casez (\$417 )
            1'h1:
                \nres_out$next  = \$422 [3:0];
          endcase
          casez (\$424 )
            1'h1:
                \nres_out$next  = \$429 [3:0];
          endcase
          casez (\$431 )
            1'h1:
                \nres_out$next  = \$436 [3:0];
          endcase
          casez (\$438 )
            1'h1:
                \nres_out$next  = \$443 [3:0];
          endcase
          casez (\$445 )
            1'h1:
                \nres_out$next  = \$450 [3:0];
          endcase
          casez (\$452 )
            1'h1:
                \nres_out$next  = \$457 [3:0];
          endcase
          casez (\$459 )
            1'h1:
                \nres_out$next  = \$464 [3:0];
          endcase
          casez (\$466 )
            1'h1:
                \nres_out$next  = \$471 [3:0];
          endcase
          casez (\$473 )
            1'h1:
                \nres_out$next  = \$478 [3:0];
          endcase
          casez (\$480 )
            1'h1:
                \nres_out$next  = \$485 [3:0];
          endcase
          casez (\$487 )
            1'h1:
                \nres_out$next  = \$492 [3:0];
          endcase
          casez (\$494 )
            1'h1:
                \nres_out$next  = \$499 [3:0];
          endcase
          casez (\$501 )
            1'h1:
                \nres_out$next  = \$506 [3:0];
          endcase
          casez (\$508 )
            1'h1:
                \nres_out$next  = \$513 [3:0];
          endcase
          casez (\$515 )
            1'h1:
                \nres_out$next  = \$520 [3:0];
          endcase
          casez (\$522 )
            1'h1:
                \nres_out$next  = \$527 [3:0];
          endcase
          casez (\$529 )
            1'h1:
                \nres_out$next  = \$534 [3:0];
          endcase
          casez (\$536 )
            1'h1:
                \nres_out$next  = \$541 [3:0];
          endcase
          casez (\$543 )
            1'h1:
                \nres_out$next  = \$548 [3:0];
          endcase
          casez (\$550 )
            1'h1:
                \nres_out$next  = \$555 [3:0];
          endcase
          casez (\$557 )
            1'h1:
                \nres_out$next  = \$562 [3:0];
          endcase
          casez (\$564 )
            1'h1:
                \nres_out$next  = \$569 [3:0];
          endcase
          casez (\$571 )
            1'h1:
                \nres_out$next  = \$576 [3:0];
          endcase
          casez (\$578 )
            1'h1:
                \nres_out$next  = \$583 [3:0];
          endcase
          casez (\$585 )
            1'h1:
                \nres_out$next  = \$590 [3:0];
          endcase
          casez (\$592 )
            1'h1:
                \nres_out$next  = \$597 [3:0];
          endcase
          casez (\$599 )
            1'h1:
                \nres_out$next  = \$604 [3:0];
          endcase
          casez (\$606 )
            1'h1:
                \nres_out$next  = \$611 [3:0];
          endcase
        end
    endcase
    casez (rst)
      1'h1:
          \nres_out$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \lastCount$next  = lastCount;
    casez (\$783 )
      1'h1:
          \lastCount$next  = t1_count;
    endcase
    casez (rst)
      1'h1:
          \lastCount$next  = 7'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    casez (\$785 )
      1'h1:
          myOutReady = 1'h0;
      default:
          myOutReady = wt_outrdy;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    bigK = 32'd0;
    casez (\$796 )
      1'h1:
          bigK = 32'd1116352408;
    endcase
    casez (\$798 )
      1'h1:
          bigK = 32'd1899447441;
    endcase
    casez (\$800 )
      1'h1:
          bigK = 32'd3049323471;
    endcase
    casez (\$802 )
      1'h1:
          bigK = 32'd3921009573;
    endcase
    casez (\$804 )
      1'h1:
          bigK = 32'd961987163;
    endcase
    casez (\$806 )
      1'h1:
          bigK = 32'd1508970993;
    endcase
    casez (\$808 )
      1'h1:
          bigK = 32'd2453635748;
    endcase
    casez (\$810 )
      1'h1:
          bigK = 32'd2870763221;
    endcase
    casez (\$812 )
      1'h1:
          bigK = 32'd3624381080;
    endcase
    casez (\$814 )
      1'h1:
          bigK = 32'd310598401;
    endcase
    casez (\$816 )
      1'h1:
          bigK = 32'd607225278;
    endcase
    casez (\$818 )
      1'h1:
          bigK = 32'd1426881987;
    endcase
    casez (\$820 )
      1'h1:
          bigK = 32'd1925078388;
    endcase
    casez (\$822 )
      1'h1:
          bigK = 32'd2162078206;
    endcase
    casez (\$824 )
      1'h1:
          bigK = 32'd2614888103;
    endcase
    casez (\$826 )
      1'h1:
          bigK = 32'd3248222580;
    endcase
    casez (\$828 )
      1'h1:
          bigK = 32'd3835390401;
    endcase
    casez (\$830 )
      1'h1:
          bigK = 32'd4022224774;
    endcase
    casez (\$832 )
      1'h1:
          bigK = 32'd264347078;
    endcase
    casez (\$834 )
      1'h1:
          bigK = 32'd604807628;
    endcase
    casez (\$836 )
      1'h1:
          bigK = 32'd770255983;
    endcase
    casez (\$838 )
      1'h1:
          bigK = 32'd1249150122;
    endcase
    casez (\$840 )
      1'h1:
          bigK = 32'd1555081692;
    endcase
    casez (\$842 )
      1'h1:
          bigK = 32'd1996064986;
    endcase
    casez (\$844 )
      1'h1:
          bigK = 32'd2554220882;
    endcase
    casez (\$846 )
      1'h1:
          bigK = 32'd2821834349;
    endcase
    casez (\$848 )
      1'h1:
          bigK = 32'd2952996808;
    endcase
    casez (\$850 )
      1'h1:
          bigK = 32'd3210313671;
    endcase
    casez (\$852 )
      1'h1:
          bigK = 32'd3336571891;
    endcase
    casez (\$854 )
      1'h1:
          bigK = 32'd3584528711;
    endcase
    casez (\$856 )
      1'h1:
          bigK = 32'd113926993;
    endcase
    casez (\$858 )
      1'h1:
          bigK = 32'd338241895;
    endcase
    casez (\$860 )
      1'h1:
          bigK = 32'd666307205;
    endcase
    casez (\$862 )
      1'h1:
          bigK = 32'd773529912;
    endcase
    casez (\$864 )
      1'h1:
          bigK = 32'd1294757372;
    endcase
    casez (\$866 )
      1'h1:
          bigK = 32'd1396182291;
    endcase
    casez (\$868 )
      1'h1:
          bigK = 32'd1695183700;
    endcase
    casez (\$870 )
      1'h1:
          bigK = 32'd1986661051;
    endcase
    casez (\$872 )
      1'h1:
          bigK = 32'd2177026350;
    endcase
    casez (\$874 )
      1'h1:
          bigK = 32'd2456956037;
    endcase
    casez (\$876 )
      1'h1:
          bigK = 32'd2730485921;
    endcase
    casez (\$878 )
      1'h1:
          bigK = 32'd2820302411;
    endcase
    casez (\$880 )
      1'h1:
          bigK = 32'd3259730800;
    endcase
    casez (\$882 )
      1'h1:
          bigK = 32'd3345764771;
    endcase
    casez (\$884 )
      1'h1:
          bigK = 32'd3516065817;
    endcase
    casez (\$886 )
      1'h1:
          bigK = 32'd3600352804;
    endcase
    casez (\$888 )
      1'h1:
          bigK = 32'd4094571909;
    endcase
    casez (\$890 )
      1'h1:
          bigK = 32'd275423344;
    endcase
    casez (\$892 )
      1'h1:
          bigK = 32'd430227734;
    endcase
    casez (\$894 )
      1'h1:
          bigK = 32'd506948616;
    endcase
    casez (\$896 )
      1'h1:
          bigK = 32'd659060556;
    endcase
    casez (\$898 )
      1'h1:
          bigK = 32'd883997877;
    endcase
    casez (\$900 )
      1'h1:
          bigK = 32'd958139571;
    endcase
    casez (\$902 )
      1'h1:
          bigK = 32'd1322822218;
    endcase
    casez (\$904 )
      1'h1:
          bigK = 32'd1537002063;
    endcase
    casez (\$906 )
      1'h1:
          bigK = 32'd1747873779;
    endcase
    casez (\$908 )
      1'h1:
          bigK = 32'd1955562222;
    endcase
    casez (\$910 )
      1'h1:
          bigK = 32'd2024104815;
    endcase
    casez (\$912 )
      1'h1:
          bigK = 32'd2227730452;
    endcase
    casez (\$914 )
      1'h1:
          bigK = 32'd2361852424;
    endcase
    casez (\$916 )
      1'h1:
          bigK = 32'd2428436474;
    endcase
    casez (\$918 )
      1'h1:
          bigK = 32'd2756734187;
    endcase
    casez (\$920 )
      1'h1:
          bigK = 32'd3204031479;
    endcase
    casez (\$922 )
      1'h1:
          bigK = 32'd3329325298;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \newMessage$next  = newMessage;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (checkedResults)
            1'h1:
                \newMessage$next  = 1'h1;
            default:
                \newMessage$next  = 1'h0;
          endcase
    endcase
    casez (rst)
      1'h1:
          \newMessage$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \wt_lastcnt$next  = wt_lastcnt;
    casez (\$931 )
      1'h1:
          \wt_lastcnt$next  = wt_count;
    endcase
    (* full_case = 32'd1 *)
    casez (\$933 )
      1'h1:
          /* empty */;
      default:
          casez (\$935 )
            1'h1:
                casez (\$937 )
                  1'h1:
                      \wt_lastcnt$next  = wt_count;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \wt_lastcnt$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \wt_outrdy$next  = wt_outrdy;
    (* full_case = 32'd1 *)
    casez (\$939 )
      1'h1:
          \wt_outrdy$next  = 1'h1;
      default:
          casez (\$941 )
            1'h1:
              begin
                casez (\$943 )
                  1'h1:
                      \wt_outrdy$next  = 1'h0;
                endcase
                casez (\$945 )
                  1'h1:
                      \wt_outrdy$next  = 1'h0;
                endcase
                casez (\$947 )
                  1'h1:
                      \wt_outrdy$next  = 1'h1;
                endcase
              end
          endcase
    endcase
    casez (rst)
      1'h1:
          \wt_outrdy$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \wt_out$next  = wt_out;
    (* full_case = 32'd1 *)
    casez (\$949 )
      1'h1:
        begin
          casez (\$951 )
            1'h1:
                \wt_out$next  = hist[511:480];
          endcase
          casez (\$953 )
            1'h1:
                \wt_out$next  = hist[479:448];
          endcase
          casez (\$955 )
            1'h1:
                \wt_out$next  = hist[447:416];
          endcase
          casez (\$957 )
            1'h1:
                \wt_out$next  = hist[415:384];
          endcase
          casez (\$959 )
            1'h1:
                \wt_out$next  = hist[383:352];
          endcase
          casez (\$961 )
            1'h1:
                \wt_out$next  = hist[351:320];
          endcase
          casez (\$963 )
            1'h1:
                \wt_out$next  = hist[319:288];
          endcase
          casez (\$965 )
            1'h1:
                \wt_out$next  = hist[287:256];
          endcase
          casez (\$967 )
            1'h1:
                \wt_out$next  = hist[255:224];
          endcase
          casez (\$969 )
            1'h1:
                \wt_out$next  = hist[223:192];
          endcase
          casez (\$971 )
            1'h1:
                \wt_out$next  = hist[191:160];
          endcase
          casez (\$973 )
            1'h1:
                \wt_out$next  = hist[159:128];
          endcase
          casez (\$975 )
            1'h1:
                \wt_out$next  = hist[127:96];
          endcase
          casez (\$977 )
            1'h1:
                \wt_out$next  = hist[95:64];
          endcase
          casez (\$979 )
            1'h1:
                \wt_out$next  = hist[63:32];
          endcase
          casez (\$981 )
            1'h1:
                \wt_out$next  = hist[31:0];
          endcase
        end
      default:
          \wt_out$next  = currentResult;
    endcase
    casez (rst)
      1'h1:
          \wt_out$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \tickDelay$next  = tickDelay;
    (* full_case = 32'd1 *)
    casez (\$983 )
      1'h1:
          /* empty */;
      default:
          casez (\$985 )
            1'h1:
              begin
                \tickDelay$next  = \$988 [1:0];
                casez (\$990 )
                  1'h1:
                      \tickDelay$next  = 2'h0;
                endcase
              end
          endcase
    endcase
    casez (rst)
      1'h1:
          \tickDelay$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \lastVal$next  = lastVal;
    (* full_case = 32'd1 *)
    casez (\$992 )
      1'h1:
          /* empty */;
      default:
          casez (\$994 )
            1'h1:
                casez (\$996 )
                  1'h1:
                      casez (\$998 )
                        1'h1:
                            \lastVal$next  = currentResult;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \lastVal$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \shiftCount$next  = shiftCount;
    (* full_case = 32'd1 *)
    casez (\$1000 )
      1'h1:
          /* empty */;
      default:
          casez (\$1002 )
            1'h1:
                casez (\$1004 )
                  1'h1:
                      casez (\$1006 )
                        1'h1:
                            \shiftCount$next  = \$1009 [8:0];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \shiftCount$next  = 9'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-1$next  = \sbuf-1 ;
    (* full_case = 32'd1 *)
    casez (\$1011 )
      1'h1:
          /* empty */;
      default:
          casez (\$1013 )
            1'h1:
                casez (\$1015 )
                  1'h1:
                      casez (\$1017 )
                        1'h1:
                            \sbuf-1$next  = hist[63:32];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-1$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in0$next  = in0;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$613 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$615 )
                        1'h1:
                            casez (\$617 )
                              1'h1:
                                  \in0$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in0$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-2$next  = \sbuf-2 ;
    (* full_case = 32'd1 *)
    casez (\$1019 )
      1'h1:
          /* empty */;
      default:
          casez (\$1021 )
            1'h1:
                casez (\$1023 )
                  1'h1:
                      casez (\$1025 )
                        1'h1:
                            \sbuf-2$next  = hist[95:64];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-2$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-3$next  = \sbuf-3 ;
    (* full_case = 32'd1 *)
    casez (\$1027 )
      1'h1:
          /* empty */;
      default:
          casez (\$1029 )
            1'h1:
                casez (\$1031 )
                  1'h1:
                      casez (\$1033 )
                        1'h1:
                            \sbuf-3$next  = hist[127:96];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-3$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-4$next  = \sbuf-4 ;
    (* full_case = 32'd1 *)
    casez (\$1035 )
      1'h1:
          /* empty */;
      default:
          casez (\$1037 )
            1'h1:
                casez (\$1039 )
                  1'h1:
                      casez (\$1041 )
                        1'h1:
                            \sbuf-4$next  = hist[159:128];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-4$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-5$next  = \sbuf-5 ;
    (* full_case = 32'd1 *)
    casez (\$1043 )
      1'h1:
          /* empty */;
      default:
          casez (\$1045 )
            1'h1:
                casez (\$1047 )
                  1'h1:
                      casez (\$1049 )
                        1'h1:
                            \sbuf-5$next  = hist[191:160];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-5$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-6$next  = \sbuf-6 ;
    (* full_case = 32'd1 *)
    casez (\$1051 )
      1'h1:
          /* empty */;
      default:
          casez (\$1053 )
            1'h1:
                casez (\$1055 )
                  1'h1:
                      casez (\$1057 )
                        1'h1:
                            \sbuf-6$next  = hist[223:192];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-6$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-7$next  = \sbuf-7 ;
    (* full_case = 32'd1 *)
    casez (\$1059 )
      1'h1:
          /* empty */;
      default:
          casez (\$1061 )
            1'h1:
                casez (\$1063 )
                  1'h1:
                      casez (\$1065 )
                        1'h1:
                            \sbuf-7$next  = hist[255:224];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-7$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-8$next  = \sbuf-8 ;
    (* full_case = 32'd1 *)
    casez (\$1067 )
      1'h1:
          /* empty */;
      default:
          casez (\$1069 )
            1'h1:
                casez (\$1071 )
                  1'h1:
                      casez (\$1073 )
                        1'h1:
                            \sbuf-8$next  = hist[287:256];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-8$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-9$next  = \sbuf-9 ;
    (* full_case = 32'd1 *)
    casez (\$1075 )
      1'h1:
          /* empty */;
      default:
          casez (\$1077 )
            1'h1:
                casez (\$1079 )
                  1'h1:
                      casez (\$1081 )
                        1'h1:
                            \sbuf-9$next  = hist[319:288];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-9$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-10$next  = \sbuf-10 ;
    (* full_case = 32'd1 *)
    casez (\$1083 )
      1'h1:
          /* empty */;
      default:
          casez (\$1085 )
            1'h1:
                casez (\$1087 )
                  1'h1:
                      casez (\$1089 )
                        1'h1:
                            \sbuf-10$next  = hist[351:320];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-10$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-11$next  = \sbuf-11 ;
    (* full_case = 32'd1 *)
    casez (\$1091 )
      1'h1:
          /* empty */;
      default:
          casez (\$1093 )
            1'h1:
                casez (\$1095 )
                  1'h1:
                      casez (\$1097 )
                        1'h1:
                            \sbuf-11$next  = hist[383:352];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-11$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in1$next  = in1;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$619 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$621 )
                        1'h1:
                            casez (\$623 )
                              1'h1:
                                  \in1$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in1$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-12$next  = \sbuf-12 ;
    (* full_case = 32'd1 *)
    casez (\$1099 )
      1'h1:
          /* empty */;
      default:
          casez (\$1101 )
            1'h1:
                casez (\$1103 )
                  1'h1:
                      casez (\$1105 )
                        1'h1:
                            \sbuf-12$next  = hist[415:384];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-12$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-13$next  = \sbuf-13 ;
    (* full_case = 32'd1 *)
    casez (\$1107 )
      1'h1:
          /* empty */;
      default:
          casez (\$1109 )
            1'h1:
                casez (\$1111 )
                  1'h1:
                      casez (\$1113 )
                        1'h1:
                            \sbuf-13$next  = hist[447:416];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-13$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-14$next  = \sbuf-14 ;
    (* full_case = 32'd1 *)
    casez (\$1115 )
      1'h1:
          /* empty */;
      default:
          casez (\$1117 )
            1'h1:
                casez (\$1119 )
                  1'h1:
                      casez (\$1121 )
                        1'h1:
                            \sbuf-14$next  = hist[479:448];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-14$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \sbuf-15$next  = \sbuf-15 ;
    (* full_case = 32'd1 *)
    casez (\$1123 )
      1'h1:
          /* empty */;
      default:
          casez (\$1125 )
            1'h1:
                casez (\$1127 )
                  1'h1:
                      casez (\$1129 )
                        1'h1:
                            \sbuf-15$next  = hist[511:480];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-15$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \debug_sig$next  = debug_sig;
    (* full_case = 32'd1 *)
    casez (\$1131 )
      1'h1:
          /* empty */;
      default:
          casez (\$1133 )
            1'h1:
                casez (\$1135 )
                  1'h1:
                      casez (\$1137 )
                        1'h1:
                            \debug_sig$next  = \$1140 [31:0];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \debug_sig$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \lastResult$next  = lastResult;
    (* full_case = 32'd1 *)
    casez (\$1142 )
      1'h1:
          /* empty */;
      default:
          casez (\$1144 )
            1'h1:
                casez (\$1146 )
                  1'h1:
                      \lastResult$next  = currentResult;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \lastResult$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \currentResult$next  = currentResult;
    (* full_case = 32'd1 *)
    casez (\$1148 )
      1'h1:
          /* empty */;
      default:
          casez (\$1150 )
            1'h1:
                casez (\$1152 )
                  1'h1:
                      \currentResult$next  = wt_res;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \currentResult$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2083:dump_module$1 ) begin end
    \in2$next  = in2;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$625 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$627 )
                        1'h1:
                            casez (\$629 )
                              1'h1:
                                  \in2$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in2$next  = 4'h0;
    endcase
  end
  assign \$1  = \$28 ;
  assign \$30  = \$31 ;
  assign \$167  = \$170 ;
  assign \$174  = \$177 ;
  assign \$181  = \$184 ;
  assign \$188  = \$191 ;
  assign \$195  = \$198 ;
  assign \$202  = \$205 ;
  assign \$209  = \$212 ;
  assign \$216  = \$219 ;
  assign \$223  = \$226 ;
  assign \$230  = \$233 ;
  assign \$237  = \$240 ;
  assign \$244  = \$247 ;
  assign \$251  = \$254 ;
  assign \$258  = \$261 ;
  assign \$265  = \$268 ;
  assign \$272  = \$275 ;
  assign \$279  = \$282 ;
  assign \$286  = \$289 ;
  assign \$293  = \$296 ;
  assign \$300  = \$303 ;
  assign \$307  = \$310 ;
  assign \$314  = \$317 ;
  assign \$321  = \$324 ;
  assign \$328  = \$331 ;
  assign \$335  = \$338 ;
  assign \$342  = \$345 ;
  assign \$349  = \$352 ;
  assign \$356  = \$359 ;
  assign \$363  = \$366 ;
  assign \$370  = \$373 ;
  assign \$377  = \$380 ;
  assign \$384  = \$387 ;
  assign \$391  = \$394 ;
  assign \$398  = \$401 ;
  assign \$405  = \$408 ;
  assign \$412  = \$415 ;
  assign \$419  = \$422 ;
  assign \$426  = \$429 ;
  assign \$433  = \$436 ;
  assign \$440  = \$443 ;
  assign \$447  = \$450 ;
  assign \$454  = \$457 ;
  assign \$461  = \$464 ;
  assign \$468  = \$471 ;
  assign \$475  = \$478 ;
  assign \$482  = \$485 ;
  assign \$489  = \$492 ;
  assign \$496  = \$499 ;
  assign \$503  = \$506 ;
  assign \$510  = \$513 ;
  assign \$517  = \$520 ;
  assign \$524  = \$527 ;
  assign \$531  = \$534 ;
  assign \$538  = \$541 ;
  assign \$545  = \$548 ;
  assign \$552  = \$555 ;
  assign \$559  = \$562 ;
  assign \$566  = \$569 ;
  assign \$573  = \$576 ;
  assign \$580  = \$583 ;
  assign \$587  = \$590 ;
  assign \$594  = \$597 ;
  assign \$601  = \$604 ;
  assign \$608  = \$611 ;
  assign \$669  = \$670 ;
  assign \$678  = \$679 ;
  assign \$725  = \$728 ;
  assign \$734  = \$735 ;
  assign \$739  = \$740 ;
  assign \$742  = \$743 ;
  assign \$745  = \$746 ;
  assign \$748  = \$749 ;
  assign \$751  = \$752 ;
  assign \$754  = \$755 ;
  assign \$757  = \$758 ;
  assign \$760  = \$761 ;
  assign \$763  = \$764 ;
  assign \$770  = \$771 ;
  assign \$773  = \$774 ;
  assign \$780  = \$781 ;
  assign \$787  = \$794 ;
  assign \$924  = \$929 ;
  assign \$987  = \$988 ;
  assign \$1008  = \$1009 ;
  assign \$1139  = \$1140 ;
  assign result = 1'h0;
  assign wt_res = \$929 [31:0];
  assign s0_s0_x = hist[479:448];
  assign s1_s1_x = hist[63:32];
  assign t1_out = \$794 [31:0];
  assign ch_ch_z = t1_g;
  assign ch_ch_y = t1_f;
  assign ch_ch_x = t1_e;
  assign rot1_rot1_x = t1_e;
  assign t1_outrdy = myOutReady;
  assign wt_count = t1_count[5:0];
  assign t2_t2_c = bp_c;
  assign t2_t2_b = bp_b;
  assign t2_t2_a = bp_a;
  assign t1_h = bp_h;
  assign t1_g = bp_g;
  assign t1_f = bp_f;
  assign t1_e = bp_e;
  assign inWord = \$28 [31:0];
  assign \$2  = { 3'h0, in0, 28'h0000000 };
  assign \$4  = { 7'h00, in1, 24'h000000 };
  assign \$8  = { 11'h000, in2, 20'h00000 };
  assign \$12  = { 15'h0000, in3, 16'h0000 };
  assign \$16  = { 3'h0, in4, 12'h000 };
  assign \$20  = { 7'h00, in5, 8'h00 };
  assign \$24  = { 3'h0, in6, 4'h0 };
  assign \$170  = { 28'h0000000, \$168 [31:28] };
  assign \$177  = { 24'h000000, \$175 [31:24] };
  assign \$184  = { 20'h00000, \$182 [31:20] };
  assign \$191  = { 16'h0000, \$189 [31:16] };
  assign \$198  = { 12'h000, \$196 [31:12] };
  assign \$205  = { 8'h00, \$203 [31:8] };
  assign \$212  = { 4'h0, \$210 [31:4] };
  assign \$219  = \$217 ;
  assign \$226  = { 28'h0000000, \$224 [31:28] };
  assign \$233  = { 24'h000000, \$231 [31:24] };
  assign \$240  = { 20'h00000, \$238 [31:20] };
  assign \$247  = { 16'h0000, \$245 [31:16] };
  assign \$254  = { 12'h000, \$252 [31:12] };
  assign \$261  = { 8'h00, \$259 [31:8] };
  assign \$268  = { 4'h0, \$266 [31:4] };
  assign \$275  = \$273 ;
  assign \$282  = { 28'h0000000, \$280 [31:28] };
  assign \$289  = { 24'h000000, \$287 [31:24] };
  assign \$296  = { 20'h00000, \$294 [31:20] };
  assign \$303  = { 16'h0000, \$301 [31:16] };
  assign \$310  = { 12'h000, \$308 [31:12] };
  assign \$317  = { 8'h00, \$315 [31:8] };
  assign \$324  = { 4'h0, \$322 [31:4] };
  assign \$331  = \$329 ;
  assign \$338  = { 28'h0000000, \$336 [31:28] };
  assign \$345  = { 24'h000000, \$343 [31:24] };
  assign \$352  = { 20'h00000, \$350 [31:20] };
  assign \$359  = { 16'h0000, \$357 [31:16] };
  assign \$366  = { 12'h000, \$364 [31:12] };
  assign \$373  = { 8'h00, \$371 [31:8] };
  assign \$380  = { 4'h0, \$378 [31:4] };
  assign \$387  = \$385 ;
  assign \$394  = { 28'h0000000, \$392 [31:28] };
  assign \$401  = { 24'h000000, \$399 [31:24] };
  assign \$408  = { 20'h00000, \$406 [31:20] };
  assign \$415  = { 16'h0000, \$413 [31:16] };
  assign \$422  = { 12'h000, \$420 [31:12] };
  assign \$429  = { 8'h00, \$427 [31:8] };
  assign \$436  = { 4'h0, \$434 [31:4] };
  assign \$443  = \$441 ;
  assign \$450  = { 28'h0000000, \$448 [31:28] };
  assign \$457  = { 24'h000000, \$455 [31:24] };
  assign \$464  = { 20'h00000, \$462 [31:20] };
  assign \$471  = { 16'h0000, \$469 [31:16] };
  assign \$478  = { 12'h000, \$476 [31:12] };
  assign \$485  = { 8'h00, \$483 [31:8] };
  assign \$492  = { 4'h0, \$490 [31:4] };
  assign \$499  = \$497 ;
  assign \$506  = { 28'h0000000, \$504 [31:28] };
  assign \$513  = { 24'h000000, \$511 [31:24] };
  assign \$520  = { 20'h00000, \$518 [31:20] };
  assign \$527  = { 16'h0000, \$525 [31:16] };
  assign \$534  = { 12'h000, \$532 [31:12] };
  assign \$541  = { 8'h00, \$539 [31:8] };
  assign \$548  = { 4'h0, \$546 [31:4] };
  assign \$555  = \$553 ;
  assign \$562  = { 28'h0000000, \$560 [31:28] };
  assign \$569  = { 24'h000000, \$567 [31:24] };
  assign \$576  = { 20'h00000, \$574 [31:20] };
  assign \$583  = { 16'h0000, \$581 [31:16] };
  assign \$590  = { 12'h000, \$588 [31:12] };
  assign \$597  = { 8'h00, \$595 [31:8] };
  assign \$604  = { 4'h0, \$602 [31:4] };
  assign \$611  = \$609 ;
  assign \$726  = { 31'h00000000, hist, 32'h00000000 };
endmodule

module psychogenic_shaman(io_in, io_out);
  wire deadPin0;
  wire deadPin1;
  wire deadPin2;
  input [7:0] io_in;
  wire [7:0] io_in;
  output [7:0] io_out;
  wire [7:0] io_out;
  wire nibbler_busy;
  wire nibbler_clk;
  wire [3:0] nibbler_inNibble;
  wire nibbler_inputReady;
  wire [3:0] nibbler_nres_out;
  wire nibbler_rst;
  nibbler nibbler (
    .busy(nibbler_busy),
    .clk(nibbler_clk),
    .inNibble(nibbler_inNibble),
    .inputReady(nibbler_inputReady),
    .nres_out(nibbler_nres_out),
    .rst(nibbler_rst)
  );
  assign io_out = { deadPin0, deadPin0, deadPin0, nibbler_busy, nibbler_nres_out };
  assign deadPin2 = 1'h0;
  assign deadPin1 = 1'h0;
  assign deadPin0 = 1'h0;
  assign nibbler_inputReady = io_in[3];
  assign nibbler_inNibble = io_in[7:4];
  assign nibbler_rst = io_in[1];
  assign nibbler_clk = io_in[0];
endmodule

module rot0(rot0_out, rot0_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] a;
  wire [31:0] b;
  wire [31:0] c;
  output [31:0] rot0_out;
  wire [31:0] rot0_out;
  input [31:0] rot0_x;
  wire [31:0] rot0_x;
  assign \$1  = a ^ b;
  assign \$3  = \$1  ^ c;
  assign rot0_out = \$3 ;
  assign c = { rot0_x[21:0], rot0_x[31:22] };
  assign b = { rot0_x[12:0], rot0_x[31:13] };
  assign a = { rot0_x[1:0], rot0_x[31:2] };
endmodule

module rot1(rot1_out, rot1_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] a;
  wire [31:0] b;
  wire [31:0] c;
  output [31:0] rot1_out;
  wire [31:0] rot1_out;
  input [31:0] rot1_x;
  wire [31:0] rot1_x;
  assign \$1  = a ^ b;
  assign \$3  = \$1  ^ c;
  assign rot1_out = \$3 ;
  assign c = { rot1_x[24:0], rot1_x[31:25] };
  assign b = { rot1_x[10:0], rot1_x[31:11] };
  assign a = { rot1_x[5:0], rot1_x[31:6] };
endmodule

module s0(s0_out, s0_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  wire [31:0] a;
  wire [31:0] b;
  wire [31:0] c;
  output [31:0] s0_out;
  wire [31:0] s0_out;
  input [31:0] s0_x;
  wire [31:0] s0_x;
  assign \$3  = a ^ b;
  assign \$5  = \$3  ^ c;
  assign s0_out = \$5 ;
  assign c = \$1 ;
  assign b = { s0_x[17:0], s0_x[31:18] };
  assign a = { s0_x[6:0], s0_x[31:7] };
  assign \$1  = { 3'h0, s0_x[31:3] };
endmodule

module s1(s1_out, s1_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  output [31:0] s1_out;
  wire [31:0] s1_out;
  input [31:0] s1_x;
  wire [31:0] s1_x;
  assign \$1  = { s1_x[16:0], s1_x[31:17] } ^ { s1_x[18:0], s1_x[31:19] };
  assign \$5  = \$1  ^ \$3 ;
  assign s1_out = \$5 ;
  assign \$3  = { 10'h000, s1_x[31:10] };
endmodule

module t2(t2_b, t2_c, t2_out, t2_a);
  wire [32:0] \$1 ;
  wire [32:0] \$2 ;
  wire [31:0] maj_maj_out;
  wire [31:0] maj_maj_x;
  wire [31:0] maj_maj_y;
  wire [31:0] maj_maj_z;
  wire [31:0] rot0_rot0_out;
  wire [31:0] rot0_rot0_x;
  input [31:0] t2_a;
  wire [31:0] t2_a;
  input [31:0] t2_b;
  wire [31:0] t2_b;
  input [31:0] t2_c;
  wire [31:0] t2_c;
  output [31:0] t2_out;
  wire [31:0] t2_out;
  assign \$2  = rot0_rot0_out + maj_maj_out;
  maj maj (
    .maj_out(maj_maj_out),
    .maj_x(maj_maj_x),
    .maj_y(maj_maj_y),
    .maj_z(maj_maj_z)
  );
  rot0 rot0 (
    .rot0_out(rot0_rot0_out),
    .rot0_x(rot0_rot0_x)
  );
  assign \$1  = \$2 ;
  assign t2_out = \$2 [31:0];
  assign maj_maj_z = t2_c;
  assign maj_maj_y = t2_b;
  assign maj_maj_x = t2_a;
  assign rot0_rot0_x = t2_a;
endmodule

