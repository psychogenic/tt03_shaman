/*
    Shama v1.0.1, for tinytapeout3.
    Copyright (C) 2023 Pat Deegan, https://psychogenic.com
    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.
    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.
    You should have received a copy of the GNU General Public License
    along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/
`default_nettype none
`timescale 1ns/1ps
/* Generated by Yosys 0.28+1 (git sha1 a9c792dce, clang 10.0.0-4ubuntu1 -fPIC -Os) */

module \buf ();
  wire \$empty_module_filler ;
endmodule

module ch(ch_y, ch_z, ch_out, ch_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  wire [31:0] \$7 ;
  output [31:0] ch_out;
  wire [31:0] ch_out;
  input [31:0] ch_x;
  wire [31:0] ch_x;
  input [31:0] ch_y;
  wire [31:0] ch_y;
  input [31:0] ch_z;
  wire [31:0] ch_z;
  assign \$1  = ch_x & ch_y;
  assign \$3  = ~ ch_x;
  assign \$5  = \$3  & ch_z;
  assign \$7  = \$1  ^ \$5 ;
  assign ch_out = \$7 ;
endmodule

module maj(maj_y, maj_z, maj_out, maj_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  wire [31:0] \$7 ;
  wire [31:0] \$9 ;
  output [31:0] maj_out;
  wire [31:0] maj_out;
  input [31:0] maj_x;
  wire [31:0] maj_x;
  input [31:0] maj_y;
  wire [31:0] maj_y;
  input [31:0] maj_z;
  wire [31:0] maj_z;
  assign \$9  = \$5  ^ \$7 ;
  assign \$1  = maj_x & maj_y;
  assign \$3  = maj_x & maj_z;
  assign \$5  = \$1  ^ \$3 ;
  assign \$7  = maj_y & maj_z;
  assign maj_out = \$9 ;
endmodule

module nibbler(rst, inNibble, inputReady, result, nres_out, busy, clk);
  reg \$auto$verilog_backend.cc:2097:dump_module$1  = 0;
  wire [34:0] \$1 ;
  wire [34:0] \$10 ;
  wire [31:0] \$100 ;
  wire \$1001 ;
  wire \$1003 ;
  wire \$1005 ;
  wire \$1007 ;
  wire \$1009 ;
  wire \$1011 ;
  wire [32:0] \$1013 ;
  wire [32:0] \$1014 ;
  wire \$1016 ;
  wire \$1018 ;
  wire \$102 ;
  wire \$1020 ;
  wire \$1022 ;
  wire \$1024 ;
  wire \$1026 ;
  wire [31:0] \$104 ;
  wire [31:0] \$105 ;
  wire [31:0] \$107 ;
  wire \$109 ;
  wire [31:0] \$111 ;
  wire [31:0] \$112 ;
  wire [31:0] \$114 ;
  wire \$116 ;
  wire [31:0] \$118 ;
  wire [31:0] \$119 ;
  wire [34:0] \$12 ;
  wire [31:0] \$121 ;
  wire \$123 ;
  wire [31:0] \$125 ;
  wire [31:0] \$126 ;
  wire [31:0] \$128 ;
  wire \$130 ;
  wire [31:0] \$132 ;
  wire [31:0] \$133 ;
  wire [31:0] \$135 ;
  wire \$137 ;
  wire [31:0] \$139 ;
  wire [34:0] \$14 ;
  wire [31:0] \$140 ;
  wire [31:0] \$142 ;
  wire \$144 ;
  wire [31:0] \$146 ;
  wire [31:0] \$147 ;
  wire [31:0] \$149 ;
  wire \$151 ;
  wire [31:0] \$153 ;
  wire [31:0] \$154 ;
  wire [31:0] \$156 ;
  wire \$158 ;
  wire [18:0] \$16 ;
  wire [31:0] \$160 ;
  wire [31:0] \$161 ;
  wire [31:0] \$163 ;
  wire \$165 ;
  wire [31:0] \$167 ;
  wire [31:0] \$168 ;
  wire [31:0] \$170 ;
  wire \$172 ;
  wire [31:0] \$174 ;
  wire [31:0] \$175 ;
  wire [31:0] \$177 ;
  wire \$179 ;
  wire [34:0] \$18 ;
  wire [31:0] \$181 ;
  wire [31:0] \$182 ;
  wire [31:0] \$184 ;
  wire \$186 ;
  wire [31:0] \$188 ;
  wire [31:0] \$189 ;
  wire [31:0] \$191 ;
  wire \$193 ;
  wire [31:0] \$195 ;
  wire [31:0] \$196 ;
  wire [31:0] \$198 ;
  wire [34:0] \$2 ;
  wire [18:0] \$20 ;
  wire \$200 ;
  wire [31:0] \$202 ;
  wire [31:0] \$203 ;
  wire [31:0] \$205 ;
  wire \$207 ;
  wire [31:0] \$209 ;
  wire [31:0] \$210 ;
  wire [31:0] \$212 ;
  wire \$214 ;
  wire [31:0] \$216 ;
  wire [31:0] \$217 ;
  wire [31:0] \$219 ;
  wire [34:0] \$22 ;
  wire \$221 ;
  wire [31:0] \$223 ;
  wire [31:0] \$224 ;
  wire [31:0] \$226 ;
  wire \$228 ;
  wire [31:0] \$230 ;
  wire [31:0] \$231 ;
  wire [31:0] \$233 ;
  wire \$235 ;
  wire [31:0] \$237 ;
  wire [31:0] \$238 ;
  wire [10:0] \$24 ;
  wire [31:0] \$240 ;
  wire \$242 ;
  wire [31:0] \$244 ;
  wire [31:0] \$245 ;
  wire [31:0] \$247 ;
  wire \$249 ;
  wire [31:0] \$251 ;
  wire [31:0] \$252 ;
  wire [31:0] \$254 ;
  wire \$256 ;
  wire [31:0] \$258 ;
  wire [31:0] \$259 ;
  wire [34:0] \$26 ;
  wire [31:0] \$261 ;
  wire \$263 ;
  wire [31:0] \$265 ;
  wire [31:0] \$266 ;
  wire [31:0] \$268 ;
  wire \$270 ;
  wire [31:0] \$272 ;
  wire [31:0] \$273 ;
  wire [31:0] \$275 ;
  wire \$277 ;
  wire [31:0] \$279 ;
  wire [34:0] \$28 ;
  wire [31:0] \$280 ;
  wire [31:0] \$282 ;
  wire \$284 ;
  wire [31:0] \$286 ;
  wire [31:0] \$287 ;
  wire [31:0] \$289 ;
  wire \$291 ;
  wire [31:0] \$293 ;
  wire [31:0] \$294 ;
  wire [31:0] \$296 ;
  wire \$298 ;
  wire [6:0] \$30 ;
  wire [31:0] \$300 ;
  wire [31:0] \$301 ;
  wire [31:0] \$303 ;
  wire \$305 ;
  wire [31:0] \$307 ;
  wire [31:0] \$308 ;
  wire [6:0] \$31 ;
  wire [31:0] \$310 ;
  wire \$312 ;
  wire [31:0] \$314 ;
  wire [31:0] \$315 ;
  wire [31:0] \$317 ;
  wire \$319 ;
  wire [31:0] \$321 ;
  wire [31:0] \$322 ;
  wire [31:0] \$324 ;
  wire \$326 ;
  wire [31:0] \$328 ;
  wire [31:0] \$329 ;
  wire \$33 ;
  wire [31:0] \$331 ;
  wire \$333 ;
  wire [31:0] \$335 ;
  wire [31:0] \$336 ;
  wire [31:0] \$338 ;
  wire \$340 ;
  wire [31:0] \$342 ;
  wire [31:0] \$343 ;
  wire [31:0] \$345 ;
  wire \$347 ;
  wire [31:0] \$349 ;
  wire \$35 ;
  wire [31:0] \$350 ;
  wire [31:0] \$352 ;
  wire \$354 ;
  wire [31:0] \$356 ;
  wire [31:0] \$357 ;
  wire [31:0] \$359 ;
  wire \$361 ;
  wire [31:0] \$363 ;
  wire [31:0] \$364 ;
  wire [31:0] \$366 ;
  wire \$368 ;
  wire \$37 ;
  wire [31:0] \$370 ;
  wire [31:0] \$371 ;
  wire [31:0] \$373 ;
  wire \$375 ;
  wire [31:0] \$377 ;
  wire [31:0] \$378 ;
  wire [31:0] \$380 ;
  wire \$382 ;
  wire [31:0] \$384 ;
  wire [31:0] \$385 ;
  wire [31:0] \$387 ;
  wire \$389 ;
  wire \$39 ;
  wire [31:0] \$391 ;
  wire [31:0] \$392 ;
  wire [31:0] \$394 ;
  wire \$396 ;
  wire [31:0] \$398 ;
  wire [31:0] \$399 ;
  wire [34:0] \$4 ;
  wire [31:0] \$401 ;
  wire \$403 ;
  wire [31:0] \$405 ;
  wire [31:0] \$406 ;
  wire [31:0] \$408 ;
  wire [31:0] \$41 ;
  wire \$410 ;
  wire [31:0] \$412 ;
  wire [31:0] \$413 ;
  wire [31:0] \$415 ;
  wire \$417 ;
  wire [31:0] \$419 ;
  wire [31:0] \$42 ;
  wire [31:0] \$420 ;
  wire [31:0] \$422 ;
  wire \$424 ;
  wire [31:0] \$426 ;
  wire [31:0] \$427 ;
  wire [31:0] \$429 ;
  wire \$431 ;
  wire [31:0] \$433 ;
  wire [31:0] \$434 ;
  wire [31:0] \$436 ;
  wire \$438 ;
  wire [31:0] \$44 ;
  wire [31:0] \$440 ;
  wire [31:0] \$441 ;
  wire [31:0] \$443 ;
  wire \$445 ;
  wire [31:0] \$447 ;
  wire [31:0] \$448 ;
  wire [31:0] \$450 ;
  wire \$452 ;
  wire [31:0] \$454 ;
  wire [31:0] \$455 ;
  wire [31:0] \$457 ;
  wire \$459 ;
  wire \$46 ;
  wire [31:0] \$461 ;
  wire [31:0] \$462 ;
  wire [31:0] \$464 ;
  wire \$466 ;
  wire [31:0] \$468 ;
  wire [31:0] \$469 ;
  wire [31:0] \$471 ;
  wire \$473 ;
  wire [31:0] \$475 ;
  wire [31:0] \$476 ;
  wire [31:0] \$478 ;
  wire [31:0] \$48 ;
  wire \$480 ;
  wire [31:0] \$482 ;
  wire [31:0] \$483 ;
  wire [31:0] \$485 ;
  wire \$487 ;
  wire \$489 ;
  wire [31:0] \$49 ;
  wire \$491 ;
  wire \$493 ;
  wire \$495 ;
  wire \$497 ;
  wire \$499 ;
  wire \$501 ;
  wire \$503 ;
  wire \$505 ;
  wire \$507 ;
  wire \$509 ;
  wire [31:0] \$51 ;
  wire \$511 ;
  wire \$513 ;
  wire \$515 ;
  wire \$517 ;
  wire \$519 ;
  wire \$521 ;
  wire \$523 ;
  wire \$525 ;
  wire \$527 ;
  wire \$529 ;
  wire \$53 ;
  wire \$531 ;
  wire \$533 ;
  wire \$535 ;
  wire \$537 ;
  wire \$539 ;
  wire \$541 ;
  wire [4:0] \$543 ;
  wire [4:0] \$544 ;
  wire \$546 ;
  wire \$548 ;
  wire [31:0] \$55 ;
  wire \$550 ;
  wire [8:0] \$552 ;
  wire [8:0] \$553 ;
  wire \$555 ;
  wire \$557 ;
  wire \$559 ;
  wire [31:0] \$56 ;
  wire \$561 ;
  wire \$563 ;
  wire \$565 ;
  wire \$567 ;
  wire \$569 ;
  wire \$571 ;
  wire \$573 ;
  wire \$575 ;
  wire \$577 ;
  wire \$579 ;
  wire [31:0] \$58 ;
  wire \$581 ;
  wire \$583 ;
  wire \$585 ;
  wire \$587 ;
  wire \$589 ;
  wire \$591 ;
  wire \$593 ;
  wire \$595 ;
  wire \$597 ;
  wire [574:0] \$599 ;
  wire [34:0] \$6 ;
  wire \$60 ;
  wire [574:0] \$600 ;
  wire [574:0] \$602 ;
  wire \$604 ;
  wire \$606 ;
  wire [5:0] \$608 ;
  wire [5:0] \$609 ;
  wire \$611 ;
  wire [7:0] \$613 ;
  wire [7:0] \$614 ;
  wire [32:0] \$616 ;
  wire [32:0] \$617 ;
  wire [32:0] \$619 ;
  wire [31:0] \$62 ;
  wire [32:0] \$620 ;
  wire [32:0] \$622 ;
  wire [32:0] \$623 ;
  wire [32:0] \$625 ;
  wire [32:0] \$626 ;
  wire [32:0] \$628 ;
  wire [32:0] \$629 ;
  wire [31:0] \$63 ;
  wire [32:0] \$631 ;
  wire [32:0] \$632 ;
  wire [32:0] \$634 ;
  wire [32:0] \$635 ;
  wire [32:0] \$637 ;
  wire [32:0] \$638 ;
  wire \$640 ;
  wire \$642 ;
  wire [32:0] \$644 ;
  wire [32:0] \$645 ;
  wire [32:0] \$647 ;
  wire [32:0] \$648 ;
  wire [31:0] \$65 ;
  wire \$650 ;
  wire \$652 ;
  wire [4:0] \$654 ;
  wire [4:0] \$655 ;
  wire \$657 ;
  wire \$659 ;
  wire [35:0] \$661 ;
  wire [32:0] \$662 ;
  wire [33:0] \$664 ;
  wire [34:0] \$666 ;
  wire [35:0] \$668 ;
  wire \$67 ;
  wire \$670 ;
  wire \$672 ;
  wire \$674 ;
  wire \$676 ;
  wire \$678 ;
  wire \$680 ;
  wire \$682 ;
  wire \$684 ;
  wire \$686 ;
  wire \$688 ;
  wire [31:0] \$69 ;
  wire \$690 ;
  wire \$692 ;
  wire \$694 ;
  wire \$696 ;
  wire \$698 ;
  wire [31:0] \$70 ;
  wire \$700 ;
  wire \$702 ;
  wire \$704 ;
  wire \$706 ;
  wire \$708 ;
  wire \$710 ;
  wire \$712 ;
  wire \$714 ;
  wire \$716 ;
  wire \$718 ;
  wire [31:0] \$72 ;
  wire \$720 ;
  wire \$722 ;
  wire \$724 ;
  wire \$726 ;
  wire \$728 ;
  wire \$730 ;
  wire \$732 ;
  wire \$734 ;
  wire \$736 ;
  wire \$738 ;
  wire \$74 ;
  wire \$740 ;
  wire \$742 ;
  wire \$744 ;
  wire \$746 ;
  wire \$748 ;
  wire \$750 ;
  wire \$752 ;
  wire \$754 ;
  wire \$756 ;
  wire \$758 ;
  wire [31:0] \$76 ;
  wire \$760 ;
  wire \$762 ;
  wire \$764 ;
  wire \$766 ;
  wire \$768 ;
  wire [31:0] \$77 ;
  wire \$770 ;
  wire \$772 ;
  wire \$774 ;
  wire \$776 ;
  wire \$778 ;
  wire \$780 ;
  wire \$782 ;
  wire \$784 ;
  wire \$786 ;
  wire \$788 ;
  wire [31:0] \$79 ;
  wire \$790 ;
  wire \$792 ;
  wire \$794 ;
  wire \$796 ;
  wire [34:0] \$798 ;
  wire [32:0] \$799 ;
  wire [34:0] \$8 ;
  wire [33:0] \$801 ;
  wire [34:0] \$803 ;
  wire \$805 ;
  wire \$807 ;
  wire \$809 ;
  wire \$81 ;
  wire \$811 ;
  wire \$813 ;
  wire \$815 ;
  wire \$817 ;
  wire \$819 ;
  wire \$821 ;
  wire \$823 ;
  wire \$825 ;
  wire \$827 ;
  wire \$829 ;
  wire [31:0] \$83 ;
  wire \$831 ;
  wire \$833 ;
  wire \$835 ;
  wire \$837 ;
  wire \$839 ;
  wire [31:0] \$84 ;
  wire \$841 ;
  wire \$843 ;
  wire \$845 ;
  wire \$847 ;
  wire \$849 ;
  wire \$851 ;
  wire \$853 ;
  wire \$855 ;
  wire \$857 ;
  wire \$859 ;
  wire [31:0] \$86 ;
  wire [2:0] \$861 ;
  wire [2:0] \$862 ;
  wire \$864 ;
  wire \$866 ;
  wire \$868 ;
  wire \$870 ;
  wire \$872 ;
  wire \$874 ;
  wire \$876 ;
  wire \$878 ;
  wire \$88 ;
  wire \$880 ;
  wire [9:0] \$882 ;
  wire [9:0] \$883 ;
  wire \$885 ;
  wire \$887 ;
  wire \$889 ;
  wire \$891 ;
  wire \$893 ;
  wire \$895 ;
  wire \$897 ;
  wire \$899 ;
  wire [31:0] \$90 ;
  wire \$901 ;
  wire \$903 ;
  wire \$905 ;
  wire \$907 ;
  wire \$909 ;
  wire [31:0] \$91 ;
  wire \$911 ;
  wire \$913 ;
  wire \$915 ;
  wire \$917 ;
  wire \$919 ;
  wire \$921 ;
  wire \$923 ;
  wire \$925 ;
  wire \$927 ;
  wire \$929 ;
  wire [31:0] \$93 ;
  wire \$931 ;
  wire \$933 ;
  wire \$935 ;
  wire \$937 ;
  wire \$939 ;
  wire \$941 ;
  wire \$943 ;
  wire \$945 ;
  wire \$947 ;
  wire \$949 ;
  wire \$95 ;
  wire \$951 ;
  wire \$953 ;
  wire \$955 ;
  wire \$957 ;
  wire \$959 ;
  wire \$961 ;
  wire \$963 ;
  wire \$965 ;
  wire \$967 ;
  wire \$969 ;
  wire [31:0] \$97 ;
  wire \$971 ;
  wire \$973 ;
  wire \$975 ;
  wire \$977 ;
  wire \$979 ;
  wire [31:0] \$98 ;
  wire \$981 ;
  wire \$983 ;
  wire \$985 ;
  wire \$987 ;
  wire \$989 ;
  wire \$991 ;
  wire \$993 ;
  wire \$995 ;
  wire \$997 ;
  wire \$999 ;
  reg [31:0] bigK;
  reg [31:0] bp_a = 32'd0;
  reg [31:0] \bp_a$next ;
  reg [31:0] bp_b = 32'd0;
  reg [31:0] \bp_b$next ;
  reg [31:0] bp_c = 32'd0;
  reg [31:0] \bp_c$next ;
  reg [31:0] bp_d = 32'd0;
  reg [31:0] \bp_d$next ;
  reg [31:0] bp_e = 32'd0;
  reg [31:0] \bp_e$next ;
  reg [31:0] bp_f = 32'd0;
  reg [31:0] \bp_f$next ;
  reg [31:0] bp_g = 32'd0;
  reg [31:0] \bp_g$next ;
  reg [31:0] bp_h = 32'd0;
  reg [31:0] \bp_h$next ;
  reg bp_outrdy = 1'h0;
  reg \bp_outrdy$next ;
  (* enum_base_type = "BlockProcessorState" *)
  (* enum_value_0000 = "PowerUp" *)
  (* enum_value_0001 = "NewMessageBegin" *)
  (* enum_value_0010 = "NewBlockBegin" *)
  (* enum_value_0011 = "WaitForReady" *)
  (* enum_value_0100 = "ValueSnapShot" *)
  (* enum_value_0101 = "ProcessBlockUnit" *)
  (* enum_value_0110 = "CheckBlockDone" *)
  (* enum_value_0111 = "ProcessBlockDone" *)
  (* enum_value_1000 = "HashReady" *)
  reg [3:0] bp_procst = 4'h0;
  reg [3:0] \bp_procst$next ;
  output busy;
  reg busy = 1'h0;
  reg \busy$next ;
  wire [31:0] ch_ch_out;
  wire [31:0] ch_ch_x;
  wire [31:0] ch_ch_y;
  wire [31:0] ch_ch_z;
  reg checkedResults = 1'h0;
  reg \checkedResults$next ;
  input clk;
  wire clk;
  reg [31:0] currentResult = 32'd0;
  reg [31:0] \currentResult$next ;
  reg [31:0] debug_sig = 32'd0;
  reg [31:0] \debug_sig$next ;
  reg [3:0] delayCount = 4'h0;
  reg [3:0] \delayCount$next ;
  reg doProcessBlock = 1'h0;
  reg \doProcessBlock$next ;
  reg [31:0] hbuf0 = 32'd0;
  reg [31:0] \hbuf0$next ;
  reg [31:0] hbuf1 = 32'd0;
  reg [31:0] \hbuf1$next ;
  reg [31:0] hbuf2 = 32'd0;
  reg [31:0] \hbuf2$next ;
  reg [31:0] hbuf3 = 32'd0;
  reg [31:0] \hbuf3$next ;
  reg [31:0] hbuf4 = 32'd0;
  reg [31:0] \hbuf4$next ;
  reg [31:0] hbuf5 = 32'd0;
  reg [31:0] \hbuf5$next ;
  reg [31:0] hbuf6 = 32'd0;
  reg [31:0] \hbuf6$next ;
  reg [31:0] hbuf7 = 32'd0;
  reg [31:0] \hbuf7$next ;
  reg [511:0] hist = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  reg [511:0] \hist$next ;
  reg [3:0] in0 = 4'h0;
  reg [3:0] \in0$next ;
  reg [3:0] in1 = 4'h0;
  reg [3:0] \in1$next ;
  reg [3:0] in2 = 4'h0;
  reg [3:0] \in2$next ;
  reg [3:0] in3 = 4'h0;
  reg [3:0] \in3$next ;
  reg [3:0] in4 = 4'h0;
  reg [3:0] \in4$next ;
  reg [3:0] in5 = 4'h0;
  reg [3:0] \in5$next ;
  reg [3:0] in6 = 4'h0;
  reg [3:0] \in6$next ;
  reg [3:0] in7 = 4'h0;
  reg [3:0] \in7$next ;
  input [3:0] inNibble;
  wire [3:0] inNibble;
  wire [31:0] inWord;
  input inputReady;
  wire inputReady;
  reg inputSeen = 1'h0;
  reg \inputSeen$next ;
  reg [6:0] lastCount = 7'h00;
  reg [6:0] \lastCount$next ;
  reg [31:0] lastResult = 32'd0;
  reg [31:0] \lastResult$next ;
  reg [31:0] lastVal = 32'd0;
  reg [31:0] \lastVal$next ;
  reg myOutReady;
  reg newMessage = 1'h0;
  reg \newMessage$next ;
  reg [7:0] nibbleCount = 8'h00;
  reg [7:0] \nibbleCount$next ;
  reg [3:0] nibbleShift = 4'h0;
  reg [3:0] \nibbleShift$next ;
  output [3:0] nres_out;
  reg [3:0] nres_out = 4'h0;
  reg [3:0] \nres_out$next ;
  reg [31:0] opT1Output = 32'd0;
  reg [31:0] \opT1Output$next ;
  reg [31:0] opT2Output = 32'd0;
  reg [31:0] \opT2Output$next ;
  input result;
  wire result;
  reg [5:0] resultOutputNibble = 6'h00;
  reg [5:0] \resultOutputNibble$next ;
  wire [31:0] rot1_rot1_out;
  wire [31:0] rot1_rot1_x;
  input rst;
  wire rst;
  wire [31:0] s0_s0_out;
  wire [31:0] s0_s0_x;
  wire [31:0] s1_s1_out;
  wire [31:0] s1_s1_x;
  reg [31:0] \sbuf-1  = 32'd0;
  reg [31:0] \sbuf-1$next ;
  reg [31:0] \sbuf-10  = 32'd0;
  reg [31:0] \sbuf-10$next ;
  reg [31:0] \sbuf-11  = 32'd0;
  reg [31:0] \sbuf-11$next ;
  reg [31:0] \sbuf-12  = 32'd0;
  reg [31:0] \sbuf-12$next ;
  reg [31:0] \sbuf-13  = 32'd0;
  reg [31:0] \sbuf-13$next ;
  reg [31:0] \sbuf-14  = 32'd0;
  reg [31:0] \sbuf-14$next ;
  reg [31:0] \sbuf-15  = 32'd0;
  reg [31:0] \sbuf-15$next ;
  reg [31:0] \sbuf-2  = 32'd0;
  reg [31:0] \sbuf-2$next ;
  reg [31:0] \sbuf-3  = 32'd0;
  reg [31:0] \sbuf-3$next ;
  reg [31:0] \sbuf-4  = 32'd0;
  reg [31:0] \sbuf-4$next ;
  reg [31:0] \sbuf-5  = 32'd0;
  reg [31:0] \sbuf-5$next ;
  reg [31:0] \sbuf-6  = 32'd0;
  reg [31:0] \sbuf-6$next ;
  reg [31:0] \sbuf-7  = 32'd0;
  reg [31:0] \sbuf-7$next ;
  reg [31:0] \sbuf-8  = 32'd0;
  reg [31:0] \sbuf-8$next ;
  reg [31:0] \sbuf-9  = 32'd0;
  reg [31:0] \sbuf-9$next ;
  reg [8:0] shiftCount = 9'h000;
  reg [8:0] \shiftCount$next ;
  reg [6:0] t1_count = 7'h00;
  reg [6:0] \t1_count$next ;
  wire [31:0] t1_e;
  wire [31:0] t1_f;
  wire [31:0] t1_g;
  wire [31:0] t1_h;
  wire [31:0] t1_out;
  wire t1_outrdy;
  wire [31:0] t2_t2_a;
  wire [31:0] t2_t2_b;
  wire [31:0] t2_t2_c;
  wire [31:0] t2_t2_out;
  reg thisIsLastUnitInBlock = 1'h0;
  reg \thisIsLastUnitInBlock$next ;
  reg [1:0] tickDelay = 2'h0;
  reg [1:0] \tickDelay$next ;
  reg [4:0] wordCount = 5'h00;
  reg [4:0] \wordCount$next ;
  wire [5:0] wt_count;
  reg [5:0] wt_lastcnt = 6'h00;
  reg [5:0] \wt_lastcnt$next ;
  reg [31:0] wt_out = 32'd0;
  reg [31:0] \wt_out$next ;
  reg wt_outrdy = 1'h0;
  reg \wt_outrdy$next ;
  wire [31:0] wt_res;
  assign \$999  = wt_count > wt_lastcnt;
  assign \$1001  = ! tickDelay;
  assign \$1003  = wt_count > 5'h10;
  assign \$1005  = wt_count < 5'h10;
  assign \$1007  = wt_count > wt_lastcnt;
  assign \$1009  = ! tickDelay;
  assign \$1011  = wt_count > 5'h10;
  assign \$1014  = debug_sig + 1'h1;
  assign \$1016  = wt_count < 5'h10;
  assign \$1018  = wt_count > wt_lastcnt;
  assign \$1020  = tickDelay == 1'h1;
  assign \$1022  = wt_count < 5'h10;
  assign \$1024  = wt_count > wt_lastcnt;
  assign \$1026  = tickDelay == 1'h1;
  always @(posedge clk)
    resultOutputNibble <= \resultOutputNibble$next ;
  always @(posedge clk)
    doProcessBlock <= \doProcessBlock$next ;
  assign \$102  = resultOutputNibble == 4'h9;
  always @(posedge clk)
    busy <= \busy$next ;
  always @(posedge clk)
    checkedResults <= \checkedResults$next ;
  always @(posedge clk)
    nres_out <= \nres_out$next ;
  always @(posedge clk)
    newMessage <= \newMessage$next ;
  always @(posedge clk)
    in0 <= \in0$next ;
  always @(posedge clk)
    in1 <= \in1$next ;
  always @(posedge clk)
    in2 <= \in2$next ;
  always @(posedge clk)
    in3 <= \in3$next ;
  always @(posedge clk)
    in4 <= \in4$next ;
  always @(posedge clk)
    in5 <= \in5$next ;
  always @(posedge clk)
    in6 <= \in6$next ;
  always @(posedge clk)
    in7 <= \in7$next ;
  always @(posedge clk)
    inputSeen <= \inputSeen$next ;
  always @(posedge clk)
    nibbleShift <= \nibbleShift$next ;
  always @(posedge clk)
    nibbleCount <= \nibbleCount$next ;
  always @(posedge clk)
    hist <= \hist$next ;
  always @(posedge clk)
    wordCount <= \wordCount$next ;
  always @(posedge clk)
    bp_procst <= \bp_procst$next ;
  always @(posedge clk)
    t1_count <= \t1_count$next ;
  always @(posedge clk)
    hbuf0 <= \hbuf0$next ;
  always @(posedge clk)
    hbuf1 <= \hbuf1$next ;
  always @(posedge clk)
    hbuf2 <= \hbuf2$next ;
  always @(posedge clk)
    hbuf3 <= \hbuf3$next ;
  always @(posedge clk)
    hbuf4 <= \hbuf4$next ;
  always @(posedge clk)
    hbuf5 <= \hbuf5$next ;
  always @(posedge clk)
    hbuf6 <= \hbuf6$next ;
  always @(posedge clk)
    hbuf7 <= \hbuf7$next ;
  always @(posedge clk)
    thisIsLastUnitInBlock <= \thisIsLastUnitInBlock$next ;
  always @(posedge clk)
    bp_outrdy <= \bp_outrdy$next ;
  always @(posedge clk)
    bp_a <= \bp_a$next ;
  always @(posedge clk)
    bp_b <= \bp_b$next ;
  always @(posedge clk)
    bp_c <= \bp_c$next ;
  always @(posedge clk)
    bp_d <= \bp_d$next ;
  always @(posedge clk)
    bp_e <= \bp_e$next ;
  always @(posedge clk)
    bp_f <= \bp_f$next ;
  always @(posedge clk)
    bp_g <= \bp_g$next ;
  always @(posedge clk)
    bp_h <= \bp_h$next ;
  always @(posedge clk)
    opT1Output <= \opT1Output$next ;
  always @(posedge clk)
    opT2Output <= \opT2Output$next ;
  always @(posedge clk)
    delayCount <= \delayCount$next ;
  always @(posedge clk)
    lastCount <= \lastCount$next ;
  always @(posedge clk)
    wt_lastcnt <= \wt_lastcnt$next ;
  always @(posedge clk)
    wt_outrdy <= \wt_outrdy$next ;
  always @(posedge clk)
    wt_out <= \wt_out$next ;
  always @(posedge clk)
    tickDelay <= \tickDelay$next ;
  always @(posedge clk)
    lastVal <= \lastVal$next ;
  always @(posedge clk)
    shiftCount <= \shiftCount$next ;
  always @(posedge clk)
    \sbuf-1  <= \sbuf-1$next ;
  always @(posedge clk)
    \sbuf-2  <= \sbuf-2$next ;
  always @(posedge clk)
    \sbuf-3  <= \sbuf-3$next ;
  always @(posedge clk)
    \sbuf-4  <= \sbuf-4$next ;
  always @(posedge clk)
    \sbuf-5  <= \sbuf-5$next ;
  always @(posedge clk)
    \sbuf-6  <= \sbuf-6$next ;
  always @(posedge clk)
    \sbuf-7  <= \sbuf-7$next ;
  always @(posedge clk)
    \sbuf-8  <= \sbuf-8$next ;
  always @(posedge clk)
    \sbuf-9  <= \sbuf-9$next ;
  always @(posedge clk)
    \sbuf-10  <= \sbuf-10$next ;
  always @(posedge clk)
    \sbuf-11  <= \sbuf-11$next ;
  always @(posedge clk)
    \sbuf-12  <= \sbuf-12$next ;
  always @(posedge clk)
    \sbuf-13  <= \sbuf-13$next ;
  always @(posedge clk)
    \sbuf-14  <= \sbuf-14$next ;
  always @(posedge clk)
    \sbuf-15  <= \sbuf-15$next ;
  always @(posedge clk)
    debug_sig <= \debug_sig$next ;
  always @(posedge clk)
    lastResult <= \lastResult$next ;
  always @(posedge clk)
    currentResult <= \currentResult$next ;
  assign \$10  = \$6  | \$8 ;
  assign \$109  = resultOutputNibble == 4'ha;
  assign \$116  = resultOutputNibble == 4'hb;
  assign \$123  = resultOutputNibble == 4'hc;
  assign \$130  = resultOutputNibble == 4'hd;
  assign \$137  = resultOutputNibble == 4'he;
  assign \$144  = resultOutputNibble == 4'hf;
  assign \$14  = \$10  | \$12 ;
  assign \$151  = resultOutputNibble == 5'h10;
  assign \$158  = resultOutputNibble == 5'h11;
  assign \$165  = resultOutputNibble == 5'h12;
  assign \$172  = resultOutputNibble == 5'h13;
  assign \$179  = resultOutputNibble == 5'h14;
  assign \$186  = resultOutputNibble == 5'h15;
  assign \$18  = \$14  | \$16 ;
  assign \$193  = resultOutputNibble == 5'h16;
  assign \$200  = resultOutputNibble == 5'h17;
  assign \$207  = resultOutputNibble == 5'h18;
  assign \$214  = resultOutputNibble == 5'h19;
  assign \$221  = resultOutputNibble == 5'h1a;
  assign \$228  = resultOutputNibble == 5'h1b;
  assign \$22  = \$18  | \$20 ;
  assign \$235  = resultOutputNibble == 5'h1c;
  assign \$242  = resultOutputNibble == 5'h1d;
  assign \$249  = resultOutputNibble == 5'h1e;
  assign \$256  = resultOutputNibble == 5'h1f;
  assign \$263  = resultOutputNibble == 6'h20;
  assign \$26  = \$22  | \$24 ;
  assign \$270  = resultOutputNibble == 6'h21;
  assign \$277  = resultOutputNibble == 6'h22;
  assign \$284  = resultOutputNibble == 6'h23;
  assign \$28  = \$26  | in7;
  assign \$291  = resultOutputNibble == 6'h24;
  assign \$298  = resultOutputNibble == 6'h25;
  assign \$305  = resultOutputNibble == 6'h26;
  assign \$312  = resultOutputNibble == 6'h27;
  assign \$31  = resultOutputNibble + 1'h1;
  assign \$319  = resultOutputNibble == 6'h28;
  assign \$326  = resultOutputNibble == 6'h29;
  assign \$333  = resultOutputNibble == 6'h2a;
  assign \$33  = nibbleCount < 8'h80;
  assign \$340  = resultOutputNibble == 6'h2b;
  assign \$347  = resultOutputNibble == 6'h2c;
  assign \$354  = resultOutputNibble == 6'h2d;
  assign \$35  = ~ busy;
  assign \$361  = resultOutputNibble == 6'h2e;
  assign \$368  = resultOutputNibble == 6'h2f;
  assign \$375  = resultOutputNibble == 6'h30;
  assign \$37  = nibbleCount < 8'h80;
  assign \$382  = resultOutputNibble == 6'h31;
  assign \$389  = resultOutputNibble == 6'h32;
  assign \$396  = resultOutputNibble == 6'h33;
  assign \$39  = ! resultOutputNibble;
  assign \$403  = resultOutputNibble == 6'h34;
  assign \$410  = resultOutputNibble == 6'h35;
  assign \$417  = resultOutputNibble == 6'h36;
  assign \$424  = resultOutputNibble == 6'h37;
  assign \$431  = resultOutputNibble == 6'h38;
  assign \$438  = resultOutputNibble == 6'h39;
  assign \$445  = resultOutputNibble == 6'h3a;
  assign \$452  = resultOutputNibble == 6'h3b;
  assign \$459  = resultOutputNibble == 6'h3c;
  assign \$466  = resultOutputNibble == 6'h3d;
  assign \$46  = resultOutputNibble == 1'h1;
  assign \$473  = resultOutputNibble == 6'h3e;
  assign \$480  = resultOutputNibble == 6'h3f;
  assign \$487  = nibbleCount < 8'h80;
  assign \$489  = ~ inputSeen;
  assign \$491  = ! nibbleShift;
  assign \$493  = nibbleCount < 8'h80;
  assign \$495  = ~ inputSeen;
  assign \$497  = nibbleShift == 1'h1;
  assign \$499  = nibbleCount < 8'h80;
  assign \$501  = ~ inputSeen;
  assign \$503  = nibbleShift == 2'h2;
  assign \$505  = nibbleCount < 8'h80;
  assign \$507  = ~ inputSeen;
  assign \$509  = nibbleShift == 2'h3;
  assign \$511  = nibbleCount < 8'h80;
  assign \$513  = ~ inputSeen;
  assign \$515  = nibbleShift == 3'h4;
  assign \$517  = nibbleCount < 8'h80;
  assign \$519  = ~ inputSeen;
  assign \$521  = nibbleShift == 3'h5;
  assign \$523  = nibbleCount < 8'h80;
  assign \$525  = ~ inputSeen;
  assign \$527  = nibbleShift == 3'h6;
  assign \$529  = nibbleCount < 8'h80;
  assign \$531  = ~ inputSeen;
  assign \$533  = nibbleShift == 3'h7;
  assign \$535  = nibbleCount < 8'h80;
  assign \$537  = ~ inputSeen;
  assign \$53  = resultOutputNibble == 2'h2;
  assign \$539  = nibbleCount < 8'h80;
  assign \$541  = ~ inputSeen;
  assign \$544  = nibbleShift + 1'h1;
  assign \$546  = nibbleShift == 4'h8;
  assign \$548  = nibbleCount < 8'h80;
  assign \$550  = ~ inputSeen;
  assign \$553  = nibbleCount + 1'h1;
  assign \$555  = nibbleCount < 8'h80;
  assign \$557  = nibbleShift == 4'h8;
  assign \$559  = ! wordCount;
  assign \$561  = wordCount == 1'h1;
  assign \$563  = wordCount == 2'h2;
  assign \$565  = wordCount == 2'h3;
  assign \$567  = wordCount == 3'h4;
  assign \$569  = wordCount == 3'h5;
  assign \$571  = wordCount == 3'h6;
  assign \$573  = wordCount == 3'h7;
  assign \$575  = wordCount == 4'h8;
  assign \$577  = wordCount == 4'h9;
  assign \$579  = wordCount == 4'ha;
  assign \$581  = wordCount == 4'hb;
  assign \$583  = wordCount == 4'hc;
  assign \$585  = wordCount == 4'hd;
  assign \$587  = wordCount == 4'he;
  assign \$589  = wordCount == 4'hf;
  assign \$591  = wt_count < 5'h10;
  assign \$593  = wt_count > wt_lastcnt;
  assign \$595  = ! tickDelay;
  assign \$597  = wt_count > 5'h10;
  assign \$602  = \$600  | currentResult;
  assign \$604  = nibbleCount < 8'h80;
  assign \$606  = nibbleShift == 4'h8;
  assign \$60  = resultOutputNibble == 2'h3;
  assign \$609  = wordCount + 1'h1;
  assign \$611  = ~ doProcessBlock;
  assign \$614  = t1_count + 1'h1;
  assign \$617  = hbuf0 + bp_a;
  assign \$620  = hbuf1 + bp_b;
  assign \$623  = hbuf2 + bp_c;
  assign \$626  = hbuf3 + bp_d;
  assign \$629  = hbuf4 + bp_e;
  assign \$632  = hbuf5 + bp_f;
  assign \$635  = hbuf6 + bp_g;
  assign \$638  = hbuf7 + bp_h;
  assign \$640  = t1_count == 6'h3f;
  assign \$642  = ~ doProcessBlock;
  assign \$645  = opT1Output + opT2Output;
  assign \$648  = bp_d + opT1Output;
  assign \$650  = lastCount != t1_count;
  assign \$652  = delayCount < 3'h4;
  assign \$655  = delayCount + 1'h1;
  assign \$657  = lastCount != t1_count;
  assign \$659  = delayCount < 3'h4;
  assign \$662  = t1_h + rot1_rot1_out;
  assign \$664  = \$662  + ch_ch_out;
  assign \$666  = \$664  + bigK;
  assign \$668  = \$666  + wt_out;
  assign \$670  = ! t1_count;
  assign \$672  = t1_count == 1'h1;
  assign \$674  = t1_count == 2'h2;
  assign \$676  = t1_count == 2'h3;
  assign \$678  = t1_count == 3'h4;
  assign \$67  = resultOutputNibble == 3'h4;
  assign \$680  = t1_count == 3'h5;
  assign \$682  = t1_count == 3'h6;
  assign \$684  = t1_count == 3'h7;
  assign \$686  = t1_count == 4'h8;
  assign \$688  = t1_count == 4'h9;
  assign \$690  = t1_count == 4'ha;
  assign \$692  = t1_count == 4'hb;
  assign \$694  = t1_count == 4'hc;
  assign \$696  = t1_count == 4'hd;
  assign \$698  = t1_count == 4'he;
  assign \$6  = \$2  | \$4 ;
  assign \$700  = t1_count == 4'hf;
  assign \$702  = t1_count == 5'h10;
  assign \$704  = t1_count == 5'h11;
  assign \$706  = t1_count == 5'h12;
  assign \$708  = t1_count == 5'h13;
  assign \$710  = t1_count == 5'h14;
  assign \$712  = t1_count == 5'h15;
  assign \$714  = t1_count == 5'h16;
  assign \$716  = t1_count == 5'h17;
  assign \$718  = t1_count == 5'h18;
  assign \$720  = t1_count == 5'h19;
  assign \$722  = t1_count == 5'h1a;
  assign \$724  = t1_count == 5'h1b;
  assign \$726  = t1_count == 5'h1c;
  assign \$728  = t1_count == 5'h1d;
  assign \$730  = t1_count == 5'h1e;
  assign \$732  = t1_count == 5'h1f;
  assign \$734  = t1_count == 6'h20;
  assign \$736  = t1_count == 6'h21;
  assign \$738  = t1_count == 6'h22;
  assign \$740  = t1_count == 6'h23;
  assign \$742  = t1_count == 6'h24;
  assign \$744  = t1_count == 6'h25;
  assign \$746  = t1_count == 6'h26;
  assign \$748  = t1_count == 6'h27;
  assign \$74  = resultOutputNibble == 3'h5;
  assign \$750  = t1_count == 6'h28;
  assign \$752  = t1_count == 6'h29;
  assign \$754  = t1_count == 6'h2a;
  assign \$756  = t1_count == 6'h2b;
  assign \$758  = t1_count == 6'h2c;
  assign \$760  = t1_count == 6'h2d;
  assign \$762  = t1_count == 6'h2e;
  assign \$764  = t1_count == 6'h2f;
  assign \$766  = t1_count == 6'h30;
  assign \$768  = t1_count == 6'h31;
  assign \$770  = t1_count == 6'h32;
  assign \$772  = t1_count == 6'h33;
  assign \$774  = t1_count == 6'h34;
  assign \$776  = t1_count == 6'h35;
  assign \$778  = t1_count == 6'h36;
  assign \$780  = t1_count == 6'h37;
  assign \$782  = t1_count == 6'h38;
  assign \$784  = t1_count == 6'h39;
  assign \$786  = t1_count == 6'h3a;
  assign \$788  = t1_count == 6'h3b;
  assign \$790  = t1_count == 6'h3c;
  assign \$792  = t1_count == 6'h3d;
  assign \$794  = t1_count == 6'h3e;
  assign \$796  = t1_count == 6'h3f;
  assign \$799  = s1_s1_out + hist[223:192];
  assign \$801  = \$799  + s0_s0_out;
  assign \$803  = \$801  + hist[511:480];
  assign \$805  = wt_lastcnt > wt_count;
  assign \$807  = wt_count < 5'h10;
  assign \$809  = wt_count > wt_lastcnt;
  assign \$811  = tickDelay == 2'h2;
  assign \$813  = wt_count < 5'h10;
  assign \$815  = wt_count > wt_lastcnt;
  assign \$817  = ! tickDelay;
  assign \$81  = resultOutputNibble == 3'h6;
  assign \$819  = tickDelay == 1'h1;
  assign \$821  = tickDelay == 2'h2;
  assign \$823  = wt_count < 5'h10;
  assign \$825  = ! wt_count;
  assign \$827  = wt_count == 1'h1;
  assign \$829  = wt_count == 2'h2;
  assign \$831  = wt_count == 2'h3;
  assign \$833  = wt_count == 3'h4;
  assign \$835  = wt_count == 3'h5;
  assign \$837  = wt_count == 3'h6;
  assign \$839  = wt_count == 3'h7;
  assign \$841  = wt_count == 4'h8;
  assign \$843  = wt_count == 4'h9;
  assign \$845  = wt_count == 4'ha;
  assign \$847  = wt_count == 4'hb;
  assign \$849  = wt_count == 4'hc;
  assign \$851  = wt_count == 4'hd;
  assign \$853  = wt_count == 4'he;
  assign \$855  = wt_count == 4'hf;
  assign \$857  = wt_count < 5'h10;
  assign \$859  = wt_count > wt_lastcnt;
  assign \$862  = tickDelay + 1'h1;
  assign \$864  = tickDelay == 2'h2;
  assign \$866  = wt_count < 5'h10;
  assign \$868  = wt_count > wt_lastcnt;
  assign \$870  = ! tickDelay;
  assign \$872  = wt_count > 5'h10;
  assign \$874  = wt_count < 5'h10;
  assign \$876  = wt_count > wt_lastcnt;
  assign \$878  = ! tickDelay;
  assign \$880  = wt_count > 5'h10;
  assign \$883  = shiftCount + 1'h1;
  assign \$885  = wt_count < 5'h10;
  assign \$887  = wt_count > wt_lastcnt;
  assign \$88  = resultOutputNibble == 3'h7;
  assign \$889  = ! tickDelay;
  assign \$891  = wt_count > 5'h10;
  assign \$893  = wt_count < 5'h10;
  assign \$895  = wt_count > wt_lastcnt;
  assign \$897  = ! tickDelay;
  assign \$899  = wt_count > 5'h10;
  assign \$901  = wt_count < 5'h10;
  assign \$903  = wt_count > wt_lastcnt;
  assign \$905  = ! tickDelay;
  assign \$907  = wt_count > 5'h10;
  assign \$909  = wt_count < 5'h10;
  assign \$911  = wt_count > wt_lastcnt;
  assign \$913  = ! tickDelay;
  assign \$915  = wt_count > 5'h10;
  assign \$917  = wt_count < 5'h10;
  assign \$919  = wt_count > wt_lastcnt;
  assign \$921  = ! tickDelay;
  assign \$923  = wt_count > 5'h10;
  assign \$925  = wt_count < 5'h10;
  assign \$927  = wt_count > wt_lastcnt;
  assign \$929  = ! tickDelay;
  assign \$931  = wt_count > 5'h10;
  assign \$933  = wt_count < 5'h10;
  assign \$935  = wt_count > wt_lastcnt;
  assign \$937  = ! tickDelay;
  assign \$939  = wt_count > 5'h10;
  assign \$941  = wt_count < 5'h10;
  assign \$943  = wt_count > wt_lastcnt;
  assign \$945  = ! tickDelay;
  assign \$947  = wt_count > 5'h10;
  assign \$949  = wt_count < 5'h10;
  assign \$951  = wt_count > wt_lastcnt;
  assign \$953  = ! tickDelay;
  assign \$955  = wt_count > 5'h10;
  assign \$957  = wt_count < 5'h10;
  assign \$95  = resultOutputNibble == 4'h8;
  assign \$959  = wt_count > wt_lastcnt;
  assign \$961  = ! tickDelay;
  assign \$963  = wt_count > 5'h10;
  assign \$965  = wt_count < 5'h10;
  assign \$967  = wt_count > wt_lastcnt;
  assign \$969  = ! tickDelay;
  assign \$971  = wt_count > 5'h10;
  assign \$973  = wt_count < 5'h10;
  assign \$975  = wt_count > wt_lastcnt;
  assign \$977  = ! tickDelay;
  assign \$979  = wt_count > 5'h10;
  assign \$981  = wt_count < 5'h10;
  assign \$983  = wt_count > wt_lastcnt;
  assign \$985  = ! tickDelay;
  assign \$987  = wt_count > 5'h10;
  assign \$989  = wt_count < 5'h10;
  assign \$991  = wt_count > wt_lastcnt;
  assign \$993  = ! tickDelay;
  assign \$995  = wt_count > 5'h10;
  assign \$997  = wt_count < 5'h10;
  \buf  \buf  (
  );
  ch ch (
    .ch_out(ch_ch_out),
    .ch_x(ch_ch_x),
    .ch_y(ch_ch_y),
    .ch_z(ch_ch_z)
  );
  rot1 rot1 (
    .rot1_out(rot1_rot1_out),
    .rot1_x(rot1_rot1_x)
  );
  s0 s0 (
    .s0_out(s0_s0_out),
    .s0_x(s0_s0_x)
  );
  s1 s1 (
    .s1_out(s1_s1_out),
    .s1_x(s1_s1_x)
  );
  t2 t2 (
    .t2_a(t2_t2_a),
    .t2_b(t2_t2_b),
    .t2_c(t2_t2_c),
    .t2_out(t2_t2_out)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \resultOutputNibble$next  = resultOutputNibble;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          \resultOutputNibble$next  = \$31 [5:0];
      default:
          casez (checkedResults)
            1'h1:
                \resultOutputNibble$next  = 6'h00;
          endcase
    endcase
    casez (rst)
      1'h1:
          \resultOutputNibble$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in3$next  = in3;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$505 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$507 )
                        1'h1:
                            casez (\$509 )
                              1'h1:
                                  \in3$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in3$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in4$next  = in4;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$511 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$513 )
                        1'h1:
                            casez (\$515 )
                              1'h1:
                                  \in4$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in4$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in5$next  = in5;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$517 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$519 )
                        1'h1:
                            casez (\$521 )
                              1'h1:
                                  \in5$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in5$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in6$next  = in6;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$523 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$525 )
                        1'h1:
                            casez (\$527 )
                              1'h1:
                                  \in6$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in6$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in7$next  = in7;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$529 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$531 )
                        1'h1:
                            casez (\$533 )
                              1'h1:
                                  \in7$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in7$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \inputSeen$next  = inputSeen;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$535 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      casez (\$537 )
                        1'h1:
                            \inputSeen$next  = 1'h1;
                      endcase
                  default:
                      \inputSeen$next  = 1'h0;
                endcase
            default:
                casez (inputSeen)
                  1'h1:
                      \inputSeen$next  = 1'h0;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \inputSeen$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \nibbleShift$next  = nibbleShift;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$539 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      casez (\$541 )
                        1'h1:
                            \nibbleShift$next  = \$544 [3:0];
                      endcase
                  default:
                      casez (\$546 )
                        1'h1:
                            casez (inputSeen)
                              1'h1:
                                  \nibbleShift$next  = 4'h0;
                            endcase
                      endcase
                endcase
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      /* empty */;
                  default:
                      casez (bp_outrdy)
                        1'h1:
                            \nibbleShift$next  = 4'h0;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \nibbleShift$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \nibbleCount$next  = nibbleCount;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$548 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$550 )
                        1'h1:
                            \nibbleCount$next  = \$553 [7:0];
                      endcase
                endcase
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      /* empty */;
                  default:
                      casez (bp_outrdy)
                        1'h1:
                            \nibbleCount$next  = 8'h00;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \nibbleCount$next  = 8'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hist$next  = hist;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$555 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      /* empty */;
                  default:
                      casez (\$557 )
                        1'h1:
                            casez (inputSeen)
                              1'h1:
                                begin
                                  casez (\$559 )
                                    1'h1:
                                        \hist$next [511:480] = inWord;
                                  endcase
                                  casez (\$561 )
                                    1'h1:
                                        \hist$next [479:448] = inWord;
                                  endcase
                                  casez (\$563 )
                                    1'h1:
                                        \hist$next [447:416] = inWord;
                                  endcase
                                  casez (\$565 )
                                    1'h1:
                                        \hist$next [415:384] = inWord;
                                  endcase
                                  casez (\$567 )
                                    1'h1:
                                        \hist$next [383:352] = inWord;
                                  endcase
                                  casez (\$569 )
                                    1'h1:
                                        \hist$next [351:320] = inWord;
                                  endcase
                                  casez (\$571 )
                                    1'h1:
                                        \hist$next [319:288] = inWord;
                                  endcase
                                  casez (\$573 )
                                    1'h1:
                                        \hist$next [287:256] = inWord;
                                  endcase
                                  casez (\$575 )
                                    1'h1:
                                        \hist$next [255:224] = inWord;
                                  endcase
                                  casez (\$577 )
                                    1'h1:
                                        \hist$next [223:192] = inWord;
                                  endcase
                                  casez (\$579 )
                                    1'h1:
                                        \hist$next [191:160] = inWord;
                                  endcase
                                  casez (\$581 )
                                    1'h1:
                                        \hist$next [159:128] = inWord;
                                  endcase
                                  casez (\$583 )
                                    1'h1:
                                        \hist$next [127:96] = inWord;
                                  endcase
                                  casez (\$585 )
                                    1'h1:
                                        \hist$next [95:64] = inWord;
                                  endcase
                                  casez (\$587 )
                                    1'h1:
                                        \hist$next [63:32] = inWord;
                                  endcase
                                  casez (\$589 )
                                    1'h1:
                                        \hist$next [31:0] = inWord;
                                  endcase
                                end
                            endcase
                      endcase
                endcase
            default:
                casez (inputSeen)
                  1'h1:
                      \hist$next [31:0] = inWord;
                endcase
          endcase
    endcase
    (* full_case = 32'd1 *)
    casez (\$591 )
      1'h1:
          /* empty */;
      default:
          casez (\$593 )
            1'h1:
                casez (\$595 )
                  1'h1:
                      casez (\$597 )
                        1'h1:
                            \hist$next  = \$602 [511:0];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \hist$next  = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \wordCount$next  = wordCount;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (\$604 )
            1'h1:
                (* full_case = 32'd1 *)
                casez (inputReady)
                  1'h1:
                      /* empty */;
                  default:
                      casez (\$606 )
                        1'h1:
                            casez (inputSeen)
                              1'h1:
                                  \wordCount$next  = \$609 [4:0];
                            endcase
                      endcase
                endcase
            default:
                casez (inputSeen)
                  1'h1:
                      \wordCount$next  = 5'h00;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \wordCount$next  = 5'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \doProcessBlock$next  = doProcessBlock;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          \doProcessBlock$next  = 1'h0;
      default:
          (* full_case = 32'd1 *)
          casez (\$33 )
            1'h1:
                \doProcessBlock$next  = 1'h0;
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      /* empty */;
                  default:
                      \doProcessBlock$next  = 1'h1;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \doProcessBlock$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_procst$next  = bp_procst;
    (* full_case = 32'd1 *)
    casez (bp_procst)
      4'h0:
          \bp_procst$next  = 4'h1;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \bp_procst$next  = 4'h2;
          endcase
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_procst$next  = 4'h3;
          endcase
      4'h3:
          casez (t1_outrdy)
            1'h1:
                \bp_procst$next  = 4'h4;
          endcase
      4'h4:
          \bp_procst$next  = 4'h5;
      4'h5:
          \bp_procst$next  = 4'h6;
      4'h6:
          (* full_case = 32'd1 *)
          casez (thisIsLastUnitInBlock)
            1'h1:
                \bp_procst$next  = 4'h7;
            default:
                \bp_procst$next  = 4'h3;
          endcase
      4'h7:
          \bp_procst$next  = 4'h8;
      4'h8:
          casez (\$611 )
            1'h1:
                \bp_procst$next  = 4'h2;
          endcase
      default:
          \bp_procst$next  = 4'h0;
    endcase
    casez (newMessage)
      1'h1:
          \bp_procst$next  = 4'h0;
    endcase
    casez (rst)
      1'h1:
          \bp_procst$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \t1_count$next  = t1_count;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \t1_count$next  = 7'h00;
          endcase
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \t1_count$next  = 7'h00;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \t1_count$next  = \$614 [6:0];
    endcase
    casez (rst)
      1'h1:
          \t1_count$next  = 7'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf0$next  = hbuf0;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf0$next  = 32'd1779033703;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf0$next  = \$617 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf0$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          \busy$next  = \$35 ;
      default:
          (* full_case = 32'd1 *)
          casez (\$37 )
            1'h1:
                \busy$next  = 1'h0;
            default:
                (* full_case = 32'd1 *)
                casez (inputSeen)
                  1'h1:
                      \busy$next  = 1'h1;
                  default:
                      (* full_case = 32'd1 *)
                      casez (bp_outrdy)
                        1'h1:
                            \busy$next  = 1'h0;
                        default:
                            \busy$next  = 1'h1;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \busy$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf1$next  = hbuf1;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf1$next  = 32'd3144134277;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf1$next  = \$620 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf1$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf2$next  = hbuf2;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf2$next  = 32'd1013904242;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf2$next  = \$623 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf2$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf3$next  = hbuf3;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf3$next  = 32'd2773480762;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf3$next  = \$626 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf3$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf4$next  = hbuf4;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf4$next  = 32'd1359893119;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf4$next  = \$629 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf4$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf5$next  = hbuf5;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf5$next  = 32'd2600822924;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf5$next  = \$632 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf5$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf6$next  = hbuf6;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf6$next  = 32'd528734635;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf6$next  = \$635 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf6$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \hbuf7$next  = hbuf7;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          casez (doProcessBlock)
            1'h1:
                \hbuf7$next  = 32'd1541459225;
          endcase
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          \hbuf7$next  = \$638 [31:0];
    endcase
    casez (rst)
      1'h1:
          \hbuf7$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \thisIsLastUnitInBlock$next  = thisIsLastUnitInBlock;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \thisIsLastUnitInBlock$next  = 1'h0;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          casez (\$640 )
            1'h1:
                \thisIsLastUnitInBlock$next  = 1'h1;
          endcase
    endcase
    casez (rst)
      1'h1:
          \thisIsLastUnitInBlock$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_outrdy$next  = bp_outrdy;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_outrdy$next  = 1'h0;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          /* empty */;
      4'h6:
          /* empty */;
      4'h7:
          /* empty */;
      4'h8:
        begin
          \bp_outrdy$next  = 1'h1;
          casez (\$642 )
            1'h1:
                \bp_outrdy$next  = 1'h0;
          endcase
        end
    endcase
    casez (rst)
      1'h1:
          \bp_outrdy$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_a$next  = bp_a;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_a$next  = hbuf0;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_a$next  = \$645 [31:0];
    endcase
    casez (rst)
      1'h1:
          \bp_a$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \checkedResults$next  = checkedResults;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          \checkedResults$next  = 1'h1;
      default:
          casez (checkedResults)
            1'h1:
                \checkedResults$next  = 1'h0;
          endcase
    endcase
    casez (rst)
      1'h1:
          \checkedResults$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_b$next  = bp_b;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_b$next  = hbuf1;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_b$next  = bp_a;
    endcase
    casez (rst)
      1'h1:
          \bp_b$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_c$next  = bp_c;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_c$next  = hbuf2;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_c$next  = bp_b;
    endcase
    casez (rst)
      1'h1:
          \bp_c$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_d$next  = bp_d;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_d$next  = hbuf3;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_d$next  = bp_c;
    endcase
    casez (rst)
      1'h1:
          \bp_d$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_e$next  = bp_e;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_e$next  = hbuf4;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_e$next  = \$648 [31:0];
    endcase
    casez (rst)
      1'h1:
          \bp_e$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_f$next  = bp_f;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_f$next  = hbuf5;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_f$next  = bp_e;
    endcase
    casez (rst)
      1'h1:
          \bp_f$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_g$next  = bp_g;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_g$next  = hbuf6;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_g$next  = bp_f;
    endcase
    casez (rst)
      1'h1:
          \bp_g$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \bp_h$next  = bp_h;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          casez (doProcessBlock)
            1'h1:
                \bp_h$next  = hbuf7;
          endcase
      4'h3:
          /* empty */;
      4'h4:
          /* empty */;
      4'h5:
          \bp_h$next  = bp_g;
    endcase
    casez (rst)
      1'h1:
          \bp_h$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \opT1Output$next  = opT1Output;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          \opT1Output$next  = t1_out;
    endcase
    casez (rst)
      1'h1:
          \opT1Output$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \opT2Output$next  = opT2Output;
    casez (bp_procst)
      4'h0:
          /* empty */;
      4'h1:
          /* empty */;
      4'h2:
          /* empty */;
      4'h3:
          /* empty */;
      4'h4:
          \opT2Output$next  = t2_t2_out;
    endcase
    casez (rst)
      1'h1:
          \opT2Output$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \delayCount$next  = delayCount;
    casez (\$650 )
      1'h1:
          \delayCount$next  = 4'h0;
    endcase
    casez (\$652 )
      1'h1:
          \delayCount$next  = \$655 [3:0];
    endcase
    casez (rst)
      1'h1:
          \delayCount$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \nres_out$next  = nres_out;
    casez (result)
      1'h1:
        begin
          casez (\$39 )
            1'h1:
                \nres_out$next  = \$44 [3:0];
          endcase
          casez (\$46 )
            1'h1:
                \nres_out$next  = \$51 [3:0];
          endcase
          casez (\$53 )
            1'h1:
                \nres_out$next  = \$58 [3:0];
          endcase
          casez (\$60 )
            1'h1:
                \nres_out$next  = \$65 [3:0];
          endcase
          casez (\$67 )
            1'h1:
                \nres_out$next  = \$72 [3:0];
          endcase
          casez (\$74 )
            1'h1:
                \nres_out$next  = \$79 [3:0];
          endcase
          casez (\$81 )
            1'h1:
                \nres_out$next  = \$86 [3:0];
          endcase
          casez (\$88 )
            1'h1:
                \nres_out$next  = \$93 [3:0];
          endcase
          casez (\$95 )
            1'h1:
                \nres_out$next  = \$100 [3:0];
          endcase
          casez (\$102 )
            1'h1:
                \nres_out$next  = \$107 [3:0];
          endcase
          casez (\$109 )
            1'h1:
                \nres_out$next  = \$114 [3:0];
          endcase
          casez (\$116 )
            1'h1:
                \nres_out$next  = \$121 [3:0];
          endcase
          casez (\$123 )
            1'h1:
                \nres_out$next  = \$128 [3:0];
          endcase
          casez (\$130 )
            1'h1:
                \nres_out$next  = \$135 [3:0];
          endcase
          casez (\$137 )
            1'h1:
                \nres_out$next  = \$142 [3:0];
          endcase
          casez (\$144 )
            1'h1:
                \nres_out$next  = \$149 [3:0];
          endcase
          casez (\$151 )
            1'h1:
                \nres_out$next  = \$156 [3:0];
          endcase
          casez (\$158 )
            1'h1:
                \nres_out$next  = \$163 [3:0];
          endcase
          casez (\$165 )
            1'h1:
                \nres_out$next  = \$170 [3:0];
          endcase
          casez (\$172 )
            1'h1:
                \nres_out$next  = \$177 [3:0];
          endcase
          casez (\$179 )
            1'h1:
                \nres_out$next  = \$184 [3:0];
          endcase
          casez (\$186 )
            1'h1:
                \nres_out$next  = \$191 [3:0];
          endcase
          casez (\$193 )
            1'h1:
                \nres_out$next  = \$198 [3:0];
          endcase
          casez (\$200 )
            1'h1:
                \nres_out$next  = \$205 [3:0];
          endcase
          casez (\$207 )
            1'h1:
                \nres_out$next  = \$212 [3:0];
          endcase
          casez (\$214 )
            1'h1:
                \nres_out$next  = \$219 [3:0];
          endcase
          casez (\$221 )
            1'h1:
                \nres_out$next  = \$226 [3:0];
          endcase
          casez (\$228 )
            1'h1:
                \nres_out$next  = \$233 [3:0];
          endcase
          casez (\$235 )
            1'h1:
                \nres_out$next  = \$240 [3:0];
          endcase
          casez (\$242 )
            1'h1:
                \nres_out$next  = \$247 [3:0];
          endcase
          casez (\$249 )
            1'h1:
                \nres_out$next  = \$254 [3:0];
          endcase
          casez (\$256 )
            1'h1:
                \nres_out$next  = \$261 [3:0];
          endcase
          casez (\$263 )
            1'h1:
                \nres_out$next  = \$268 [3:0];
          endcase
          casez (\$270 )
            1'h1:
                \nres_out$next  = \$275 [3:0];
          endcase
          casez (\$277 )
            1'h1:
                \nres_out$next  = \$282 [3:0];
          endcase
          casez (\$284 )
            1'h1:
                \nres_out$next  = \$289 [3:0];
          endcase
          casez (\$291 )
            1'h1:
                \nres_out$next  = \$296 [3:0];
          endcase
          casez (\$298 )
            1'h1:
                \nres_out$next  = \$303 [3:0];
          endcase
          casez (\$305 )
            1'h1:
                \nres_out$next  = \$310 [3:0];
          endcase
          casez (\$312 )
            1'h1:
                \nres_out$next  = \$317 [3:0];
          endcase
          casez (\$319 )
            1'h1:
                \nres_out$next  = \$324 [3:0];
          endcase
          casez (\$326 )
            1'h1:
                \nres_out$next  = \$331 [3:0];
          endcase
          casez (\$333 )
            1'h1:
                \nres_out$next  = \$338 [3:0];
          endcase
          casez (\$340 )
            1'h1:
                \nres_out$next  = \$345 [3:0];
          endcase
          casez (\$347 )
            1'h1:
                \nres_out$next  = \$352 [3:0];
          endcase
          casez (\$354 )
            1'h1:
                \nres_out$next  = \$359 [3:0];
          endcase
          casez (\$361 )
            1'h1:
                \nres_out$next  = \$366 [3:0];
          endcase
          casez (\$368 )
            1'h1:
                \nres_out$next  = \$373 [3:0];
          endcase
          casez (\$375 )
            1'h1:
                \nres_out$next  = \$380 [3:0];
          endcase
          casez (\$382 )
            1'h1:
                \nres_out$next  = \$387 [3:0];
          endcase
          casez (\$389 )
            1'h1:
                \nres_out$next  = \$394 [3:0];
          endcase
          casez (\$396 )
            1'h1:
                \nres_out$next  = \$401 [3:0];
          endcase
          casez (\$403 )
            1'h1:
                \nres_out$next  = \$408 [3:0];
          endcase
          casez (\$410 )
            1'h1:
                \nres_out$next  = \$415 [3:0];
          endcase
          casez (\$417 )
            1'h1:
                \nres_out$next  = \$422 [3:0];
          endcase
          casez (\$424 )
            1'h1:
                \nres_out$next  = \$429 [3:0];
          endcase
          casez (\$431 )
            1'h1:
                \nres_out$next  = \$436 [3:0];
          endcase
          casez (\$438 )
            1'h1:
                \nres_out$next  = \$443 [3:0];
          endcase
          casez (\$445 )
            1'h1:
                \nres_out$next  = \$450 [3:0];
          endcase
          casez (\$452 )
            1'h1:
                \nres_out$next  = \$457 [3:0];
          endcase
          casez (\$459 )
            1'h1:
                \nres_out$next  = \$464 [3:0];
          endcase
          casez (\$466 )
            1'h1:
                \nres_out$next  = \$471 [3:0];
          endcase
          casez (\$473 )
            1'h1:
                \nres_out$next  = \$478 [3:0];
          endcase
          casez (\$480 )
            1'h1:
                \nres_out$next  = \$485 [3:0];
          endcase
        end
    endcase
    casez (rst)
      1'h1:
          \nres_out$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \lastCount$next  = lastCount;
    casez (\$657 )
      1'h1:
          \lastCount$next  = t1_count;
    endcase
    casez (rst)
      1'h1:
          \lastCount$next  = 7'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    casez (\$659 )
      1'h1:
          myOutReady = 1'h0;
      default:
          myOutReady = wt_outrdy;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    bigK = 32'd0;
    casez (\$670 )
      1'h1:
          bigK = 32'd1116352408;
    endcase
    casez (\$672 )
      1'h1:
          bigK = 32'd1899447441;
    endcase
    casez (\$674 )
      1'h1:
          bigK = 32'd3049323471;
    endcase
    casez (\$676 )
      1'h1:
          bigK = 32'd3921009573;
    endcase
    casez (\$678 )
      1'h1:
          bigK = 32'd961987163;
    endcase
    casez (\$680 )
      1'h1:
          bigK = 32'd1508970993;
    endcase
    casez (\$682 )
      1'h1:
          bigK = 32'd2453635748;
    endcase
    casez (\$684 )
      1'h1:
          bigK = 32'd2870763221;
    endcase
    casez (\$686 )
      1'h1:
          bigK = 32'd3624381080;
    endcase
    casez (\$688 )
      1'h1:
          bigK = 32'd310598401;
    endcase
    casez (\$690 )
      1'h1:
          bigK = 32'd607225278;
    endcase
    casez (\$692 )
      1'h1:
          bigK = 32'd1426881987;
    endcase
    casez (\$694 )
      1'h1:
          bigK = 32'd1925078388;
    endcase
    casez (\$696 )
      1'h1:
          bigK = 32'd2162078206;
    endcase
    casez (\$698 )
      1'h1:
          bigK = 32'd2614888103;
    endcase
    casez (\$700 )
      1'h1:
          bigK = 32'd3248222580;
    endcase
    casez (\$702 )
      1'h1:
          bigK = 32'd3835390401;
    endcase
    casez (\$704 )
      1'h1:
          bigK = 32'd4022224774;
    endcase
    casez (\$706 )
      1'h1:
          bigK = 32'd264347078;
    endcase
    casez (\$708 )
      1'h1:
          bigK = 32'd604807628;
    endcase
    casez (\$710 )
      1'h1:
          bigK = 32'd770255983;
    endcase
    casez (\$712 )
      1'h1:
          bigK = 32'd1249150122;
    endcase
    casez (\$714 )
      1'h1:
          bigK = 32'd1555081692;
    endcase
    casez (\$716 )
      1'h1:
          bigK = 32'd1996064986;
    endcase
    casez (\$718 )
      1'h1:
          bigK = 32'd2554220882;
    endcase
    casez (\$720 )
      1'h1:
          bigK = 32'd2821834349;
    endcase
    casez (\$722 )
      1'h1:
          bigK = 32'd2952996808;
    endcase
    casez (\$724 )
      1'h1:
          bigK = 32'd3210313671;
    endcase
    casez (\$726 )
      1'h1:
          bigK = 32'd3336571891;
    endcase
    casez (\$728 )
      1'h1:
          bigK = 32'd3584528711;
    endcase
    casez (\$730 )
      1'h1:
          bigK = 32'd113926993;
    endcase
    casez (\$732 )
      1'h1:
          bigK = 32'd338241895;
    endcase
    casez (\$734 )
      1'h1:
          bigK = 32'd666307205;
    endcase
    casez (\$736 )
      1'h1:
          bigK = 32'd773529912;
    endcase
    casez (\$738 )
      1'h1:
          bigK = 32'd1294757372;
    endcase
    casez (\$740 )
      1'h1:
          bigK = 32'd1396182291;
    endcase
    casez (\$742 )
      1'h1:
          bigK = 32'd1695183700;
    endcase
    casez (\$744 )
      1'h1:
          bigK = 32'd1986661051;
    endcase
    casez (\$746 )
      1'h1:
          bigK = 32'd2177026350;
    endcase
    casez (\$748 )
      1'h1:
          bigK = 32'd2456956037;
    endcase
    casez (\$750 )
      1'h1:
          bigK = 32'd2730485921;
    endcase
    casez (\$752 )
      1'h1:
          bigK = 32'd2820302411;
    endcase
    casez (\$754 )
      1'h1:
          bigK = 32'd3259730800;
    endcase
    casez (\$756 )
      1'h1:
          bigK = 32'd3345764771;
    endcase
    casez (\$758 )
      1'h1:
          bigK = 32'd3516065817;
    endcase
    casez (\$760 )
      1'h1:
          bigK = 32'd3600352804;
    endcase
    casez (\$762 )
      1'h1:
          bigK = 32'd4094571909;
    endcase
    casez (\$764 )
      1'h1:
          bigK = 32'd275423344;
    endcase
    casez (\$766 )
      1'h1:
          bigK = 32'd430227734;
    endcase
    casez (\$768 )
      1'h1:
          bigK = 32'd506948616;
    endcase
    casez (\$770 )
      1'h1:
          bigK = 32'd659060556;
    endcase
    casez (\$772 )
      1'h1:
          bigK = 32'd883997877;
    endcase
    casez (\$774 )
      1'h1:
          bigK = 32'd958139571;
    endcase
    casez (\$776 )
      1'h1:
          bigK = 32'd1322822218;
    endcase
    casez (\$778 )
      1'h1:
          bigK = 32'd1537002063;
    endcase
    casez (\$780 )
      1'h1:
          bigK = 32'd1747873779;
    endcase
    casez (\$782 )
      1'h1:
          bigK = 32'd1955562222;
    endcase
    casez (\$784 )
      1'h1:
          bigK = 32'd2024104815;
    endcase
    casez (\$786 )
      1'h1:
          bigK = 32'd2227730452;
    endcase
    casez (\$788 )
      1'h1:
          bigK = 32'd2361852424;
    endcase
    casez (\$790 )
      1'h1:
          bigK = 32'd2428436474;
    endcase
    casez (\$792 )
      1'h1:
          bigK = 32'd2756734187;
    endcase
    casez (\$794 )
      1'h1:
          bigK = 32'd3204031479;
    endcase
    casez (\$796 )
      1'h1:
          bigK = 32'd3329325298;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \newMessage$next  = newMessage;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          (* full_case = 32'd1 *)
          casez (checkedResults)
            1'h1:
                \newMessage$next  = 1'h1;
            default:
                \newMessage$next  = 1'h0;
          endcase
    endcase
    casez (rst)
      1'h1:
          \newMessage$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \wt_lastcnt$next  = wt_lastcnt;
    casez (\$805 )
      1'h1:
          \wt_lastcnt$next  = wt_count;
    endcase
    (* full_case = 32'd1 *)
    casez (\$807 )
      1'h1:
          /* empty */;
      default:
          casez (\$809 )
            1'h1:
                casez (\$811 )
                  1'h1:
                      \wt_lastcnt$next  = wt_count;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \wt_lastcnt$next  = 6'h00;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \wt_outrdy$next  = wt_outrdy;
    (* full_case = 32'd1 *)
    casez (\$813 )
      1'h1:
          \wt_outrdy$next  = 1'h1;
      default:
          casez (\$815 )
            1'h1:
              begin
                casez (\$817 )
                  1'h1:
                      \wt_outrdy$next  = 1'h0;
                endcase
                casez (\$819 )
                  1'h1:
                      \wt_outrdy$next  = 1'h0;
                endcase
                casez (\$821 )
                  1'h1:
                      \wt_outrdy$next  = 1'h1;
                endcase
              end
          endcase
    endcase
    casez (rst)
      1'h1:
          \wt_outrdy$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \wt_out$next  = wt_out;
    (* full_case = 32'd1 *)
    casez (\$823 )
      1'h1:
        begin
          casez (\$825 )
            1'h1:
                \wt_out$next  = hist[511:480];
          endcase
          casez (\$827 )
            1'h1:
                \wt_out$next  = hist[479:448];
          endcase
          casez (\$829 )
            1'h1:
                \wt_out$next  = hist[447:416];
          endcase
          casez (\$831 )
            1'h1:
                \wt_out$next  = hist[415:384];
          endcase
          casez (\$833 )
            1'h1:
                \wt_out$next  = hist[383:352];
          endcase
          casez (\$835 )
            1'h1:
                \wt_out$next  = hist[351:320];
          endcase
          casez (\$837 )
            1'h1:
                \wt_out$next  = hist[319:288];
          endcase
          casez (\$839 )
            1'h1:
                \wt_out$next  = hist[287:256];
          endcase
          casez (\$841 )
            1'h1:
                \wt_out$next  = hist[255:224];
          endcase
          casez (\$843 )
            1'h1:
                \wt_out$next  = hist[223:192];
          endcase
          casez (\$845 )
            1'h1:
                \wt_out$next  = hist[191:160];
          endcase
          casez (\$847 )
            1'h1:
                \wt_out$next  = hist[159:128];
          endcase
          casez (\$849 )
            1'h1:
                \wt_out$next  = hist[127:96];
          endcase
          casez (\$851 )
            1'h1:
                \wt_out$next  = hist[95:64];
          endcase
          casez (\$853 )
            1'h1:
                \wt_out$next  = hist[63:32];
          endcase
          casez (\$855 )
            1'h1:
                \wt_out$next  = hist[31:0];
          endcase
        end
      default:
          \wt_out$next  = currentResult;
    endcase
    casez (rst)
      1'h1:
          \wt_out$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \tickDelay$next  = tickDelay;
    (* full_case = 32'd1 *)
    casez (\$857 )
      1'h1:
          /* empty */;
      default:
          casez (\$859 )
            1'h1:
              begin
                \tickDelay$next  = \$862 [1:0];
                casez (\$864 )
                  1'h1:
                      \tickDelay$next  = 2'h0;
                endcase
              end
          endcase
    endcase
    casez (rst)
      1'h1:
          \tickDelay$next  = 2'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \lastVal$next  = lastVal;
    (* full_case = 32'd1 *)
    casez (\$866 )
      1'h1:
          /* empty */;
      default:
          casez (\$868 )
            1'h1:
                casez (\$870 )
                  1'h1:
                      casez (\$872 )
                        1'h1:
                            \lastVal$next  = currentResult;
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \lastVal$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \shiftCount$next  = shiftCount;
    (* full_case = 32'd1 *)
    casez (\$874 )
      1'h1:
          /* empty */;
      default:
          casez (\$876 )
            1'h1:
                casez (\$878 )
                  1'h1:
                      casez (\$880 )
                        1'h1:
                            \shiftCount$next  = \$883 [8:0];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \shiftCount$next  = 9'h000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-1$next  = \sbuf-1 ;
    (* full_case = 32'd1 *)
    casez (\$885 )
      1'h1:
          /* empty */;
      default:
          casez (\$887 )
            1'h1:
                casez (\$889 )
                  1'h1:
                      casez (\$891 )
                        1'h1:
                            \sbuf-1$next  = hist[63:32];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-1$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in0$next  = in0;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$487 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$489 )
                        1'h1:
                            casez (\$491 )
                              1'h1:
                                  \in0$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in0$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-2$next  = \sbuf-2 ;
    (* full_case = 32'd1 *)
    casez (\$893 )
      1'h1:
          /* empty */;
      default:
          casez (\$895 )
            1'h1:
                casez (\$897 )
                  1'h1:
                      casez (\$899 )
                        1'h1:
                            \sbuf-2$next  = hist[95:64];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-2$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-3$next  = \sbuf-3 ;
    (* full_case = 32'd1 *)
    casez (\$901 )
      1'h1:
          /* empty */;
      default:
          casez (\$903 )
            1'h1:
                casez (\$905 )
                  1'h1:
                      casez (\$907 )
                        1'h1:
                            \sbuf-3$next  = hist[127:96];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-3$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-4$next  = \sbuf-4 ;
    (* full_case = 32'd1 *)
    casez (\$909 )
      1'h1:
          /* empty */;
      default:
          casez (\$911 )
            1'h1:
                casez (\$913 )
                  1'h1:
                      casez (\$915 )
                        1'h1:
                            \sbuf-4$next  = hist[159:128];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-4$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-5$next  = \sbuf-5 ;
    (* full_case = 32'd1 *)
    casez (\$917 )
      1'h1:
          /* empty */;
      default:
          casez (\$919 )
            1'h1:
                casez (\$921 )
                  1'h1:
                      casez (\$923 )
                        1'h1:
                            \sbuf-5$next  = hist[191:160];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-5$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-6$next  = \sbuf-6 ;
    (* full_case = 32'd1 *)
    casez (\$925 )
      1'h1:
          /* empty */;
      default:
          casez (\$927 )
            1'h1:
                casez (\$929 )
                  1'h1:
                      casez (\$931 )
                        1'h1:
                            \sbuf-6$next  = hist[223:192];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-6$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-7$next  = \sbuf-7 ;
    (* full_case = 32'd1 *)
    casez (\$933 )
      1'h1:
          /* empty */;
      default:
          casez (\$935 )
            1'h1:
                casez (\$937 )
                  1'h1:
                      casez (\$939 )
                        1'h1:
                            \sbuf-7$next  = hist[255:224];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-7$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-8$next  = \sbuf-8 ;
    (* full_case = 32'd1 *)
    casez (\$941 )
      1'h1:
          /* empty */;
      default:
          casez (\$943 )
            1'h1:
                casez (\$945 )
                  1'h1:
                      casez (\$947 )
                        1'h1:
                            \sbuf-8$next  = hist[287:256];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-8$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-9$next  = \sbuf-9 ;
    (* full_case = 32'd1 *)
    casez (\$949 )
      1'h1:
          /* empty */;
      default:
          casez (\$951 )
            1'h1:
                casez (\$953 )
                  1'h1:
                      casez (\$955 )
                        1'h1:
                            \sbuf-9$next  = hist[319:288];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-9$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-10$next  = \sbuf-10 ;
    (* full_case = 32'd1 *)
    casez (\$957 )
      1'h1:
          /* empty */;
      default:
          casez (\$959 )
            1'h1:
                casez (\$961 )
                  1'h1:
                      casez (\$963 )
                        1'h1:
                            \sbuf-10$next  = hist[351:320];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-10$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-11$next  = \sbuf-11 ;
    (* full_case = 32'd1 *)
    casez (\$965 )
      1'h1:
          /* empty */;
      default:
          casez (\$967 )
            1'h1:
                casez (\$969 )
                  1'h1:
                      casez (\$971 )
                        1'h1:
                            \sbuf-11$next  = hist[383:352];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-11$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in1$next  = in1;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$493 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$495 )
                        1'h1:
                            casez (\$497 )
                              1'h1:
                                  \in1$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in1$next  = 4'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-12$next  = \sbuf-12 ;
    (* full_case = 32'd1 *)
    casez (\$973 )
      1'h1:
          /* empty */;
      default:
          casez (\$975 )
            1'h1:
                casez (\$977 )
                  1'h1:
                      casez (\$979 )
                        1'h1:
                            \sbuf-12$next  = hist[415:384];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-12$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-13$next  = \sbuf-13 ;
    (* full_case = 32'd1 *)
    casez (\$981 )
      1'h1:
          /* empty */;
      default:
          casez (\$983 )
            1'h1:
                casez (\$985 )
                  1'h1:
                      casez (\$987 )
                        1'h1:
                            \sbuf-13$next  = hist[447:416];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-13$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-14$next  = \sbuf-14 ;
    (* full_case = 32'd1 *)
    casez (\$989 )
      1'h1:
          /* empty */;
      default:
          casez (\$991 )
            1'h1:
                casez (\$993 )
                  1'h1:
                      casez (\$995 )
                        1'h1:
                            \sbuf-14$next  = hist[479:448];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-14$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \sbuf-15$next  = \sbuf-15 ;
    (* full_case = 32'd1 *)
    casez (\$997 )
      1'h1:
          /* empty */;
      default:
          casez (\$999 )
            1'h1:
                casez (\$1001 )
                  1'h1:
                      casez (\$1003 )
                        1'h1:
                            \sbuf-15$next  = hist[511:480];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \sbuf-15$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \debug_sig$next  = debug_sig;
    (* full_case = 32'd1 *)
    casez (\$1005 )
      1'h1:
          /* empty */;
      default:
          casez (\$1007 )
            1'h1:
                casez (\$1009 )
                  1'h1:
                      casez (\$1011 )
                        1'h1:
                            \debug_sig$next  = \$1014 [31:0];
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \debug_sig$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \lastResult$next  = lastResult;
    (* full_case = 32'd1 *)
    casez (\$1016 )
      1'h1:
          /* empty */;
      default:
          casez (\$1018 )
            1'h1:
                casez (\$1020 )
                  1'h1:
                      \lastResult$next  = currentResult;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \lastResult$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \currentResult$next  = currentResult;
    (* full_case = 32'd1 *)
    casez (\$1022 )
      1'h1:
          /* empty */;
      default:
          casez (\$1024 )
            1'h1:
                casez (\$1026 )
                  1'h1:
                      \currentResult$next  = wt_res;
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \currentResult$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \in2$next  = in2;
    (* full_case = 32'd1 *)
    casez (result)
      1'h1:
          /* empty */;
      default:
          casez (\$499 )
            1'h1:
                casez (inputReady)
                  1'h1:
                      casez (\$501 )
                        1'h1:
                            casez (\$503 )
                              1'h1:
                                  \in2$next  = inNibble;
                            endcase
                      endcase
                endcase
          endcase
    endcase
    casez (rst)
      1'h1:
          \in2$next  = 4'h0;
    endcase
  end
  assign \$1  = \$28 ;
  assign \$30  = \$31 ;
  assign \$41  = \$44 ;
  assign \$48  = \$51 ;
  assign \$55  = \$58 ;
  assign \$62  = \$65 ;
  assign \$69  = \$72 ;
  assign \$76  = \$79 ;
  assign \$83  = \$86 ;
  assign \$90  = \$93 ;
  assign \$97  = \$100 ;
  assign \$104  = \$107 ;
  assign \$111  = \$114 ;
  assign \$118  = \$121 ;
  assign \$125  = \$128 ;
  assign \$132  = \$135 ;
  assign \$139  = \$142 ;
  assign \$146  = \$149 ;
  assign \$153  = \$156 ;
  assign \$160  = \$163 ;
  assign \$167  = \$170 ;
  assign \$174  = \$177 ;
  assign \$181  = \$184 ;
  assign \$188  = \$191 ;
  assign \$195  = \$198 ;
  assign \$202  = \$205 ;
  assign \$209  = \$212 ;
  assign \$216  = \$219 ;
  assign \$223  = \$226 ;
  assign \$230  = \$233 ;
  assign \$237  = \$240 ;
  assign \$244  = \$247 ;
  assign \$251  = \$254 ;
  assign \$258  = \$261 ;
  assign \$265  = \$268 ;
  assign \$272  = \$275 ;
  assign \$279  = \$282 ;
  assign \$286  = \$289 ;
  assign \$293  = \$296 ;
  assign \$300  = \$303 ;
  assign \$307  = \$310 ;
  assign \$314  = \$317 ;
  assign \$321  = \$324 ;
  assign \$328  = \$331 ;
  assign \$335  = \$338 ;
  assign \$342  = \$345 ;
  assign \$349  = \$352 ;
  assign \$356  = \$359 ;
  assign \$363  = \$366 ;
  assign \$370  = \$373 ;
  assign \$377  = \$380 ;
  assign \$384  = \$387 ;
  assign \$391  = \$394 ;
  assign \$398  = \$401 ;
  assign \$405  = \$408 ;
  assign \$412  = \$415 ;
  assign \$419  = \$422 ;
  assign \$426  = \$429 ;
  assign \$433  = \$436 ;
  assign \$440  = \$443 ;
  assign \$447  = \$450 ;
  assign \$454  = \$457 ;
  assign \$461  = \$464 ;
  assign \$468  = \$471 ;
  assign \$475  = \$478 ;
  assign \$482  = \$485 ;
  assign \$543  = \$544 ;
  assign \$552  = \$553 ;
  assign \$599  = \$602 ;
  assign \$608  = \$609 ;
  assign \$613  = \$614 ;
  assign \$616  = \$617 ;
  assign \$619  = \$620 ;
  assign \$622  = \$623 ;
  assign \$625  = \$626 ;
  assign \$628  = \$629 ;
  assign \$631  = \$632 ;
  assign \$634  = \$635 ;
  assign \$637  = \$638 ;
  assign \$644  = \$645 ;
  assign \$647  = \$648 ;
  assign \$654  = \$655 ;
  assign \$661  = \$668 ;
  assign \$798  = \$803 ;
  assign \$861  = \$862 ;
  assign \$882  = \$883 ;
  assign \$1013  = \$1014 ;
  assign wt_res = \$803 [31:0];
  assign s0_s0_x = hist[479:448];
  assign s1_s1_x = hist[63:32];
  assign t1_out = \$668 [31:0];
  assign ch_ch_z = t1_g;
  assign ch_ch_y = t1_f;
  assign ch_ch_x = t1_e;
  assign rot1_rot1_x = t1_e;
  assign t1_outrdy = myOutReady;
  assign wt_count = t1_count[5:0];
  assign t2_t2_c = bp_c;
  assign t2_t2_b = bp_b;
  assign t2_t2_a = bp_a;
  assign t1_h = bp_h;
  assign t1_g = bp_g;
  assign t1_f = bp_f;
  assign t1_e = bp_e;
  assign inWord = \$28 [31:0];
  assign \$2  = { 3'h0, in0, 28'h0000000 };
  assign \$4  = { 7'h00, in1, 24'h000000 };
  assign \$8  = { 11'h000, in2, 20'h00000 };
  assign \$12  = { 15'h0000, in3, 16'h0000 };
  assign \$16  = { 3'h0, in4, 12'h000 };
  assign \$20  = { 7'h00, in5, 8'h00 };
  assign \$24  = { 3'h0, in6, 4'h0 };
  assign \$42 [27:0] = 28'h0000000;
  assign \$42 [31:28] = hbuf0[31:28];
  assign \$44  = { 28'h0000000, hbuf0[31:28] };
  assign { \$49 [31:28], \$49 [23:0] } = 28'h0000000;
  assign \$49 [27:24] = hbuf0[27:24];
  assign \$51  = { 28'h0000000, hbuf0[27:24] };
  assign { \$56 [31:24], \$56 [19:0] } = 28'h0000000;
  assign \$56 [23:20] = hbuf0[23:20];
  assign \$58  = { 28'h0000000, hbuf0[23:20] };
  assign { \$63 [31:20], \$63 [15:0] } = 28'h0000000;
  assign \$63 [19:16] = hbuf0[19:16];
  assign \$65  = { 28'h0000000, hbuf0[19:16] };
  assign { \$70 [31:16], \$70 [11:0] } = 28'h0000000;
  assign \$70 [15:12] = hbuf0[15:12];
  assign \$72  = { 28'h0000000, hbuf0[15:12] };
  assign { \$77 [31:12], \$77 [7:0] } = 28'h0000000;
  assign \$77 [11:8] = hbuf0[11:8];
  assign \$79  = { 28'h0000000, hbuf0[11:8] };
  assign { \$84 [31:8], \$84 [3:0] } = 28'h0000000;
  assign \$84 [7:4] = hbuf0[7:4];
  assign \$86  = { 28'h0000000, hbuf0[7:4] };
  assign \$91 [31:4] = 28'h0000000;
  assign \$91 [3:0] = hbuf0[3:0];
  assign \$93  = { 28'h0000000, hbuf0[3:0] };
  assign \$98 [27:0] = 28'h0000000;
  assign \$98 [31:28] = hbuf1[31:28];
  assign \$100  = { 28'h0000000, hbuf1[31:28] };
  assign { \$105 [31:28], \$105 [23:0] } = 28'h0000000;
  assign \$105 [27:24] = hbuf1[27:24];
  assign \$107  = { 28'h0000000, hbuf1[27:24] };
  assign { \$112 [31:24], \$112 [19:0] } = 28'h0000000;
  assign \$112 [23:20] = hbuf1[23:20];
  assign \$114  = { 28'h0000000, hbuf1[23:20] };
  assign { \$119 [31:20], \$119 [15:0] } = 28'h0000000;
  assign \$119 [19:16] = hbuf1[19:16];
  assign \$121  = { 28'h0000000, hbuf1[19:16] };
  assign { \$126 [31:16], \$126 [11:0] } = 28'h0000000;
  assign \$126 [15:12] = hbuf1[15:12];
  assign \$128  = { 28'h0000000, hbuf1[15:12] };
  assign { \$133 [31:12], \$133 [7:0] } = 28'h0000000;
  assign \$133 [11:8] = hbuf1[11:8];
  assign \$135  = { 28'h0000000, hbuf1[11:8] };
  assign { \$140 [31:8], \$140 [3:0] } = 28'h0000000;
  assign \$140 [7:4] = hbuf1[7:4];
  assign \$142  = { 28'h0000000, hbuf1[7:4] };
  assign \$147 [31:4] = 28'h0000000;
  assign \$147 [3:0] = hbuf1[3:0];
  assign \$149  = { 28'h0000000, hbuf1[3:0] };
  assign \$154 [27:0] = 28'h0000000;
  assign \$154 [31:28] = hbuf2[31:28];
  assign \$156  = { 28'h0000000, hbuf2[31:28] };
  assign { \$161 [31:28], \$161 [23:0] } = 28'h0000000;
  assign \$161 [27:24] = hbuf2[27:24];
  assign \$163  = { 28'h0000000, hbuf2[27:24] };
  assign { \$168 [31:24], \$168 [19:0] } = 28'h0000000;
  assign \$168 [23:20] = hbuf2[23:20];
  assign \$170  = { 28'h0000000, hbuf2[23:20] };
  assign { \$175 [31:20], \$175 [15:0] } = 28'h0000000;
  assign \$175 [19:16] = hbuf2[19:16];
  assign \$177  = { 28'h0000000, hbuf2[19:16] };
  assign { \$182 [31:16], \$182 [11:0] } = 28'h0000000;
  assign \$182 [15:12] = hbuf2[15:12];
  assign \$184  = { 28'h0000000, hbuf2[15:12] };
  assign { \$189 [31:12], \$189 [7:0] } = 28'h0000000;
  assign \$189 [11:8] = hbuf2[11:8];
  assign \$191  = { 28'h0000000, hbuf2[11:8] };
  assign { \$196 [31:8], \$196 [3:0] } = 28'h0000000;
  assign \$196 [7:4] = hbuf2[7:4];
  assign \$198  = { 28'h0000000, hbuf2[7:4] };
  assign \$203 [31:4] = 28'h0000000;
  assign \$203 [3:0] = hbuf2[3:0];
  assign \$205  = { 28'h0000000, hbuf2[3:0] };
  assign \$210 [27:0] = 28'h0000000;
  assign \$210 [31:28] = hbuf3[31:28];
  assign \$212  = { 28'h0000000, hbuf3[31:28] };
  assign { \$217 [31:28], \$217 [23:0] } = 28'h0000000;
  assign \$217 [27:24] = hbuf3[27:24];
  assign \$219  = { 28'h0000000, hbuf3[27:24] };
  assign { \$224 [31:24], \$224 [19:0] } = 28'h0000000;
  assign \$224 [23:20] = hbuf3[23:20];
  assign \$226  = { 28'h0000000, hbuf3[23:20] };
  assign { \$231 [31:20], \$231 [15:0] } = 28'h0000000;
  assign \$231 [19:16] = hbuf3[19:16];
  assign \$233  = { 28'h0000000, hbuf3[19:16] };
  assign { \$238 [31:16], \$238 [11:0] } = 28'h0000000;
  assign \$238 [15:12] = hbuf3[15:12];
  assign \$240  = { 28'h0000000, hbuf3[15:12] };
  assign { \$245 [31:12], \$245 [7:0] } = 28'h0000000;
  assign \$245 [11:8] = hbuf3[11:8];
  assign \$247  = { 28'h0000000, hbuf3[11:8] };
  assign { \$252 [31:8], \$252 [3:0] } = 28'h0000000;
  assign \$252 [7:4] = hbuf3[7:4];
  assign \$254  = { 28'h0000000, hbuf3[7:4] };
  assign \$259 [31:4] = 28'h0000000;
  assign \$259 [3:0] = hbuf3[3:0];
  assign \$261  = { 28'h0000000, hbuf3[3:0] };
  assign \$266 [27:0] = 28'h0000000;
  assign \$266 [31:28] = hbuf4[31:28];
  assign \$268  = { 28'h0000000, hbuf4[31:28] };
  assign { \$273 [31:28], \$273 [23:0] } = 28'h0000000;
  assign \$273 [27:24] = hbuf4[27:24];
  assign \$275  = { 28'h0000000, hbuf4[27:24] };
  assign { \$280 [31:24], \$280 [19:0] } = 28'h0000000;
  assign \$280 [23:20] = hbuf4[23:20];
  assign \$282  = { 28'h0000000, hbuf4[23:20] };
  assign { \$287 [31:20], \$287 [15:0] } = 28'h0000000;
  assign \$287 [19:16] = hbuf4[19:16];
  assign \$289  = { 28'h0000000, hbuf4[19:16] };
  assign { \$294 [31:16], \$294 [11:0] } = 28'h0000000;
  assign \$294 [15:12] = hbuf4[15:12];
  assign \$296  = { 28'h0000000, hbuf4[15:12] };
  assign { \$301 [31:12], \$301 [7:0] } = 28'h0000000;
  assign \$301 [11:8] = hbuf4[11:8];
  assign \$303  = { 28'h0000000, hbuf4[11:8] };
  assign { \$308 [31:8], \$308 [3:0] } = 28'h0000000;
  assign \$308 [7:4] = hbuf4[7:4];
  assign \$310  = { 28'h0000000, hbuf4[7:4] };
  assign \$315 [31:4] = 28'h0000000;
  assign \$315 [3:0] = hbuf4[3:0];
  assign \$317  = { 28'h0000000, hbuf4[3:0] };
  assign \$322 [27:0] = 28'h0000000;
  assign \$322 [31:28] = hbuf5[31:28];
  assign \$324  = { 28'h0000000, hbuf5[31:28] };
  assign { \$329 [31:28], \$329 [23:0] } = 28'h0000000;
  assign \$329 [27:24] = hbuf5[27:24];
  assign \$331  = { 28'h0000000, hbuf5[27:24] };
  assign { \$336 [31:24], \$336 [19:0] } = 28'h0000000;
  assign \$336 [23:20] = hbuf5[23:20];
  assign \$338  = { 28'h0000000, hbuf5[23:20] };
  assign { \$343 [31:20], \$343 [15:0] } = 28'h0000000;
  assign \$343 [19:16] = hbuf5[19:16];
  assign \$345  = { 28'h0000000, hbuf5[19:16] };
  assign { \$350 [31:16], \$350 [11:0] } = 28'h0000000;
  assign \$350 [15:12] = hbuf5[15:12];
  assign \$352  = { 28'h0000000, hbuf5[15:12] };
  assign { \$357 [31:12], \$357 [7:0] } = 28'h0000000;
  assign \$357 [11:8] = hbuf5[11:8];
  assign \$359  = { 28'h0000000, hbuf5[11:8] };
  assign { \$364 [31:8], \$364 [3:0] } = 28'h0000000;
  assign \$364 [7:4] = hbuf5[7:4];
  assign \$366  = { 28'h0000000, hbuf5[7:4] };
  assign \$371 [31:4] = 28'h0000000;
  assign \$371 [3:0] = hbuf5[3:0];
  assign \$373  = { 28'h0000000, hbuf5[3:0] };
  assign \$378 [27:0] = 28'h0000000;
  assign \$378 [31:28] = hbuf6[31:28];
  assign \$380  = { 28'h0000000, hbuf6[31:28] };
  assign { \$385 [31:28], \$385 [23:0] } = 28'h0000000;
  assign \$385 [27:24] = hbuf6[27:24];
  assign \$387  = { 28'h0000000, hbuf6[27:24] };
  assign { \$392 [31:24], \$392 [19:0] } = 28'h0000000;
  assign \$392 [23:20] = hbuf6[23:20];
  assign \$394  = { 28'h0000000, hbuf6[23:20] };
  assign { \$399 [31:20], \$399 [15:0] } = 28'h0000000;
  assign \$399 [19:16] = hbuf6[19:16];
  assign \$401  = { 28'h0000000, hbuf6[19:16] };
  assign { \$406 [31:16], \$406 [11:0] } = 28'h0000000;
  assign \$406 [15:12] = hbuf6[15:12];
  assign \$408  = { 28'h0000000, hbuf6[15:12] };
  assign { \$413 [31:12], \$413 [7:0] } = 28'h0000000;
  assign \$413 [11:8] = hbuf6[11:8];
  assign \$415  = { 28'h0000000, hbuf6[11:8] };
  assign { \$420 [31:8], \$420 [3:0] } = 28'h0000000;
  assign \$420 [7:4] = hbuf6[7:4];
  assign \$422  = { 28'h0000000, hbuf6[7:4] };
  assign \$427 [31:4] = 28'h0000000;
  assign \$427 [3:0] = hbuf6[3:0];
  assign \$429  = { 28'h0000000, hbuf6[3:0] };
  assign \$434 [27:0] = 28'h0000000;
  assign \$434 [31:28] = hbuf7[31:28];
  assign \$436  = { 28'h0000000, hbuf7[31:28] };
  assign { \$441 [31:28], \$441 [23:0] } = 28'h0000000;
  assign \$441 [27:24] = hbuf7[27:24];
  assign \$443  = { 28'h0000000, hbuf7[27:24] };
  assign { \$448 [31:24], \$448 [19:0] } = 28'h0000000;
  assign \$448 [23:20] = hbuf7[23:20];
  assign \$450  = { 28'h0000000, hbuf7[23:20] };
  assign { \$455 [31:20], \$455 [15:0] } = 28'h0000000;
  assign \$455 [19:16] = hbuf7[19:16];
  assign \$457  = { 28'h0000000, hbuf7[19:16] };
  assign { \$462 [31:16], \$462 [11:0] } = 28'h0000000;
  assign \$462 [15:12] = hbuf7[15:12];
  assign \$464  = { 28'h0000000, hbuf7[15:12] };
  assign { \$469 [31:12], \$469 [7:0] } = 28'h0000000;
  assign \$469 [11:8] = hbuf7[11:8];
  assign \$471  = { 28'h0000000, hbuf7[11:8] };
  assign { \$476 [31:8], \$476 [3:0] } = 28'h0000000;
  assign \$476 [7:4] = hbuf7[7:4];
  assign \$478  = { 28'h0000000, hbuf7[7:4] };
  assign \$483 [31:4] = 28'h0000000;
  assign \$483 [3:0] = hbuf7[3:0];
  assign \$485  = { 28'h0000000, hbuf7[3:0] };
  assign \$600  = { 31'h00000000, hist, 32'h00000000 };
endmodule

module psychogenic_shaman(io_in, io_out);
  wire deadPin0;
  wire deadPin1;
  wire deadPin2;
  input [7:0] io_in;
  wire [7:0] io_in;
  output [7:0] io_out;
  wire [7:0] io_out;
  wire nibbler_busy;
  wire nibbler_clk;
  wire [3:0] nibbler_inNibble;
  wire nibbler_inputReady;
  wire [3:0] nibbler_nres_out;
  wire nibbler_result;
  wire nibbler_rst;
  nibbler nibbler (
    .busy(nibbler_busy),
    .clk(nibbler_clk),
    .inNibble(nibbler_inNibble),
    .inputReady(nibbler_inputReady),
    .nres_out(nibbler_nres_out),
    .result(nibbler_result),
    .rst(nibbler_rst)
  );
  assign io_out[4] = nibbler_busy;
  assign io_out[3] = nibbler_nres_out[3];
  assign io_out[2] = nibbler_nres_out[2];
  assign io_out[1] = nibbler_nres_out[1];
  assign io_out[0] = nibbler_nres_out[0];
  assign io_out[7:5] = 3'h0;
  assign deadPin2 = 1'h0;
  assign deadPin1 = 1'h0;
  assign deadPin0 = 1'h0;
  assign nibbler_result = io_in[2];
  assign nibbler_inputReady = io_in[3];
  assign nibbler_inNibble[3] = io_in[7];
  assign nibbler_inNibble[2] = io_in[6];
  assign nibbler_inNibble[1] = io_in[5];
  assign nibbler_inNibble[0] = io_in[4];
  assign nibbler_rst = io_in[1];
  assign nibbler_clk = io_in[0];
endmodule

module rot0(rot0_out, rot0_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] a;
  wire [31:0] b;
  wire [31:0] c;
  output [31:0] rot0_out;
  wire [31:0] rot0_out;
  input [31:0] rot0_x;
  wire [31:0] rot0_x;
  assign \$1  = a ^ b;
  assign \$3  = \$1  ^ c;
  assign rot0_out = \$3 ;
  assign c = { rot0_x[21:0], rot0_x[31:22] };
  assign b = { rot0_x[12:0], rot0_x[31:13] };
  assign a = { rot0_x[1:0], rot0_x[31:2] };
endmodule

module rot1(rot1_out, rot1_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] a;
  wire [31:0] b;
  wire [31:0] c;
  output [31:0] rot1_out;
  wire [31:0] rot1_out;
  input [31:0] rot1_x;
  wire [31:0] rot1_x;
  assign \$1  = a ^ b;
  assign \$3  = \$1  ^ c;
  assign rot1_out = \$3 ;
  assign c = { rot1_x[24:0], rot1_x[31:25] };
  assign b = { rot1_x[10:0], rot1_x[31:11] };
  assign a = { rot1_x[5:0], rot1_x[31:6] };
endmodule

module s0(s0_out, s0_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  wire [31:0] a;
  wire [31:0] b;
  wire [31:0] c;
  output [31:0] s0_out;
  wire [31:0] s0_out;
  input [31:0] s0_x;
  wire [31:0] s0_x;
  assign \$3  = a ^ b;
  assign \$5  = \$3  ^ c;
  assign s0_out = \$5 ;
  assign c = \$1 ;
  assign b = { s0_x[17:0], s0_x[31:18] };
  assign a = { s0_x[6:0], s0_x[31:7] };
  assign \$1  = { 3'h0, s0_x[31:3] };
endmodule

module s1(s1_out, s1_x);
  wire [31:0] \$1 ;
  wire [31:0] \$3 ;
  wire [31:0] \$5 ;
  output [31:0] s1_out;
  wire [31:0] s1_out;
  input [31:0] s1_x;
  wire [31:0] s1_x;
  assign \$1  = { s1_x[16:0], s1_x[31:17] } ^ { s1_x[18:0], s1_x[31:19] };
  assign \$5  = \$1  ^ \$3 ;
  assign s1_out = \$5 ;
  assign \$3  = { 10'h000, s1_x[31:10] };
endmodule

module t2(t2_b, t2_c, t2_out, t2_a);
  wire [32:0] \$1 ;
  wire [32:0] \$2 ;
  wire [31:0] maj_maj_out;
  wire [31:0] maj_maj_x;
  wire [31:0] maj_maj_y;
  wire [31:0] maj_maj_z;
  wire [31:0] rot0_rot0_out;
  wire [31:0] rot0_rot0_x;
  input [31:0] t2_a;
  wire [31:0] t2_a;
  input [31:0] t2_b;
  wire [31:0] t2_b;
  input [31:0] t2_c;
  wire [31:0] t2_c;
  output [31:0] t2_out;
  wire [31:0] t2_out;
  assign \$2  = rot0_rot0_out + maj_maj_out;
  maj maj (
    .maj_out(maj_maj_out),
    .maj_x(maj_maj_x),
    .maj_y(maj_maj_y),
    .maj_z(maj_maj_z)
  );
  rot0 rot0 (
    .rot0_out(rot0_rot0_out),
    .rot0_x(rot0_rot0_x)
  );
  assign \$1  = \$2 ;
  assign t2_out = \$2 [31:0];
  assign maj_maj_z = t2_c;
  assign maj_maj_y = t2_b;
  assign maj_maj_x = t2_a;
  assign rot0_rot0_x = t2_a;
endmodule

